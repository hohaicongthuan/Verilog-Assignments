library verilog;
use verilog.vl_types.all;
entity TrafficLightController_vlg_vec_tst is
end TrafficLightController_vlg_vec_tst;
