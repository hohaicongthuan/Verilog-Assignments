library verilog;
use verilog.vl_types.all;
entity Controller_Outputs is
    generic(
        S0              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        S1              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        S2              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        S3              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        S4              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        S5              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        S6              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        S7              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        S8              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        S9              : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        S10             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        S11             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        S12             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        S13             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        S14             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        S15             : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        S16             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        S17             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        S18             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        S19             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        S20             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        S21             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        S22             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0);
        S23             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        S24             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        S25             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        S26             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        S27             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi1);
        S28             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        S29             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi0, Hi1);
        S30             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        S31             : vl_logic_vector(0 to 5) := (Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        S32             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        S33             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        S34             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        S35             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        S36             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        S37             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        S38             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        S39             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        S40             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        S41             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        S42             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        S43             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        S44             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi1, Hi0, Hi0);
        S45             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        S46             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        S47             : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi1);
        S48             : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        S49             : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        S50             : vl_logic_vector(0 to 5) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0)
    );
    port(
        CurrentState    : in     vl_logic_vector(5 downto 0);
        data_o          : out    vl_logic_vector(13 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S0 : constant is 1;
    attribute mti_svvh_generic_type of S1 : constant is 1;
    attribute mti_svvh_generic_type of S2 : constant is 1;
    attribute mti_svvh_generic_type of S3 : constant is 1;
    attribute mti_svvh_generic_type of S4 : constant is 1;
    attribute mti_svvh_generic_type of S5 : constant is 1;
    attribute mti_svvh_generic_type of S6 : constant is 1;
    attribute mti_svvh_generic_type of S7 : constant is 1;
    attribute mti_svvh_generic_type of S8 : constant is 1;
    attribute mti_svvh_generic_type of S9 : constant is 1;
    attribute mti_svvh_generic_type of S10 : constant is 1;
    attribute mti_svvh_generic_type of S11 : constant is 1;
    attribute mti_svvh_generic_type of S12 : constant is 1;
    attribute mti_svvh_generic_type of S13 : constant is 1;
    attribute mti_svvh_generic_type of S14 : constant is 1;
    attribute mti_svvh_generic_type of S15 : constant is 1;
    attribute mti_svvh_generic_type of S16 : constant is 1;
    attribute mti_svvh_generic_type of S17 : constant is 1;
    attribute mti_svvh_generic_type of S18 : constant is 1;
    attribute mti_svvh_generic_type of S19 : constant is 1;
    attribute mti_svvh_generic_type of S20 : constant is 1;
    attribute mti_svvh_generic_type of S21 : constant is 1;
    attribute mti_svvh_generic_type of S22 : constant is 1;
    attribute mti_svvh_generic_type of S23 : constant is 1;
    attribute mti_svvh_generic_type of S24 : constant is 1;
    attribute mti_svvh_generic_type of S25 : constant is 1;
    attribute mti_svvh_generic_type of S26 : constant is 1;
    attribute mti_svvh_generic_type of S27 : constant is 1;
    attribute mti_svvh_generic_type of S28 : constant is 1;
    attribute mti_svvh_generic_type of S29 : constant is 1;
    attribute mti_svvh_generic_type of S30 : constant is 1;
    attribute mti_svvh_generic_type of S31 : constant is 1;
    attribute mti_svvh_generic_type of S32 : constant is 1;
    attribute mti_svvh_generic_type of S33 : constant is 1;
    attribute mti_svvh_generic_type of S34 : constant is 1;
    attribute mti_svvh_generic_type of S35 : constant is 1;
    attribute mti_svvh_generic_type of S36 : constant is 1;
    attribute mti_svvh_generic_type of S37 : constant is 1;
    attribute mti_svvh_generic_type of S38 : constant is 1;
    attribute mti_svvh_generic_type of S39 : constant is 1;
    attribute mti_svvh_generic_type of S40 : constant is 1;
    attribute mti_svvh_generic_type of S41 : constant is 1;
    attribute mti_svvh_generic_type of S42 : constant is 1;
    attribute mti_svvh_generic_type of S43 : constant is 1;
    attribute mti_svvh_generic_type of S44 : constant is 1;
    attribute mti_svvh_generic_type of S45 : constant is 1;
    attribute mti_svvh_generic_type of S46 : constant is 1;
    attribute mti_svvh_generic_type of S47 : constant is 1;
    attribute mti_svvh_generic_type of S48 : constant is 1;
    attribute mti_svvh_generic_type of S49 : constant is 1;
    attribute mti_svvh_generic_type of S50 : constant is 1;
end Controller_Outputs;
