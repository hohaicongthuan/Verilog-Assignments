module LUT(data_i, data_o);
	input [11:0] data_i;
	output reg [22:0] data_o;
	
	always @ (data_i) begin
		case (data_i)
		12'd 0 : data_o = 23'b 00000000000000000000000 ;
		12'd 1 : data_o = 23'b 11111111110000000000010 ;
		12'd 2 : data_o = 23'b 11111111100000000001011 ;
		12'd 3 : data_o = 23'b 11111111010000000011010 ;
		12'd 4 : data_o = 23'b 11111111000000000101111 ;
		12'd 5 : data_o = 23'b 11111110110000001001010 ;
		12'd 6 : data_o = 23'b 11111110100000001101011 ;
		12'd 7 : data_o = 23'b 11111110010000010010010 ;
		12'd 8 : data_o = 23'b 11111110000000010111111 ;
		12'd 9 : data_o = 23'b 11111101110000011110010 ;
		12'd 10 : data_o = 23'b 11111101100000100101011 ;
		12'd 11 : data_o = 23'b 11111101010000101101001 ;
		12'd 12 : data_o = 23'b 11111101000000110101110 ;
		12'd 13 : data_o = 23'b 11111100110000111111000 ;
		12'd 14 : data_o = 23'b 11111100100001001001001 ;
		12'd 15 : data_o = 23'b 11111100010001010011111 ;
		12'd 16 : data_o = 23'b 11111100000001011111100 ;
		12'd 17 : data_o = 23'b 11111011110001101011110 ;
		12'd 18 : data_o = 23'b 11111011100001111000110 ;
		12'd 19 : data_o = 23'b 11111011010010000110100 ;
		12'd 20 : data_o = 23'b 11111011000010010101000 ;
		12'd 21 : data_o = 23'b 11111010110010100100010 ;
		12'd 22 : data_o = 23'b 11111010100010110100001 ;
		12'd 23 : data_o = 23'b 11111010010011000100111 ;
		12'd 24 : data_o = 23'b 11111010000011010110010 ;
		12'd 25 : data_o = 23'b 11111001110011101000011 ;
		12'd 26 : data_o = 23'b 11111001100011111011010 ;
		12'd 27 : data_o = 23'b 11111001010100001110111 ;
		12'd 28 : data_o = 23'b 11111001000100100011010 ;
		12'd 29 : data_o = 23'b 11111000110100111000011 ;
		12'd 30 : data_o = 23'b 11111000100101001110001 ;
		12'd 31 : data_o = 23'b 11111000010101100100110 ;
		12'd 32 : data_o = 23'b 11111000000101111100000 ;
		12'd 33 : data_o = 23'b 11110111110110010100000 ;
		12'd 34 : data_o = 23'b 11110111100110101100110 ;
		12'd 35 : data_o = 23'b 11110111010111000110001 ;
		12'd 36 : data_o = 23'b 11110111000111100000010 ;
		12'd 37 : data_o = 23'b 11110110110111111011010 ;
		12'd 38 : data_o = 23'b 11110110101000010110111 ;
		12'd 39 : data_o = 23'b 11110110011000110011001 ;
		12'd 40 : data_o = 23'b 11110110001001010000010 ;
		12'd 41 : data_o = 23'b 11110101111001101110000 ;
		12'd 42 : data_o = 23'b 11110101101010001100100 ;
		12'd 43 : data_o = 23'b 11110101011010101011110 ;
		12'd 44 : data_o = 23'b 11110101001011001011101 ;
		12'd 45 : data_o = 23'b 11110100111011101100011 ;
		12'd 46 : data_o = 23'b 11110100101100001101110 ;
		12'd 47 : data_o = 23'b 11110100011100101111111 ;
		12'd 48 : data_o = 23'b 11110100001101010010101 ;
		12'd 49 : data_o = 23'b 11110011111101110110001 ;
		12'd 50 : data_o = 23'b 11110011101110011010011 ;
		12'd 51 : data_o = 23'b 11110011011110111111011 ;
		12'd 52 : data_o = 23'b 11110011001111100101000 ;
		12'd 53 : data_o = 23'b 11110011000000001011011 ;
		12'd 54 : data_o = 23'b 11110010110000110010100 ;
		12'd 55 : data_o = 23'b 11110010100001011010011 ;
		12'd 56 : data_o = 23'b 11110010010010000010111 ;
		12'd 57 : data_o = 23'b 11110010000010101100001 ;
		12'd 58 : data_o = 23'b 11110001110011010110000 ;
		12'd 59 : data_o = 23'b 11110001100100000000101 ;
		12'd 60 : data_o = 23'b 11110001010100101100000 ;
		12'd 61 : data_o = 23'b 11110001000101011000001 ;
		12'd 62 : data_o = 23'b 11110000110110000100111 ;
		12'd 63 : data_o = 23'b 11110000100110110010011 ;
		12'd 64 : data_o = 23'b 11110000010111100000100 ;
		12'd 65 : data_o = 23'b 11110000001000001111100 ;
		12'd 66 : data_o = 23'b 11101111111000111111000 ;
		12'd 67 : data_o = 23'b 11101111101001101111011 ;
		12'd 68 : data_o = 23'b 11101111011010100000011 ;
		12'd 69 : data_o = 23'b 11101111001011010010000 ;
		12'd 70 : data_o = 23'b 11101110111100000100100 ;
		12'd 71 : data_o = 23'b 11101110101100110111100 ;
		12'd 72 : data_o = 23'b 11101110011101101011011 ;
		12'd 73 : data_o = 23'b 11101110001110011111111 ;
		12'd 74 : data_o = 23'b 11101101111111010101001 ;
		12'd 75 : data_o = 23'b 11101101110000001011000 ;
		12'd 76 : data_o = 23'b 11101101100001000001101 ;
		12'd 77 : data_o = 23'b 11101101010001111000111 ;
		12'd 78 : data_o = 23'b 11101101000010110000111 ;
		12'd 79 : data_o = 23'b 11101100110011101001100 ;
		12'd 80 : data_o = 23'b 11101100100100100010111 ;
		12'd 81 : data_o = 23'b 11101100010101011101000 ;
		12'd 82 : data_o = 23'b 11101100000110010111110 ;
		12'd 83 : data_o = 23'b 11101011110111010011010 ;
		12'd 84 : data_o = 23'b 11101011101000001111011 ;
		12'd 85 : data_o = 23'b 11101011011001001100010 ;
		12'd 86 : data_o = 23'b 11101011001010001001110 ;
		12'd 87 : data_o = 23'b 11101010111011001000000 ;
		12'd 88 : data_o = 23'b 11101010101100000110111 ;
		12'd 89 : data_o = 23'b 11101010011101000110100 ;
		12'd 90 : data_o = 23'b 11101010001110000110111 ;
		12'd 91 : data_o = 23'b 11101001111111000111110 ;
		12'd 92 : data_o = 23'b 11101001110000001001100 ;
		12'd 93 : data_o = 23'b 11101001100001001011111 ;
		12'd 94 : data_o = 23'b 11101001010010001110111 ;
		12'd 95 : data_o = 23'b 11101001000011010010101 ;
		12'd 96 : data_o = 23'b 11101000110100010111000 ;
		12'd 97 : data_o = 23'b 11101000100101011100001 ;
		12'd 98 : data_o = 23'b 11101000010110100001111 ;
		12'd 99 : data_o = 23'b 11101000000111101000011 ;
		12'd 100 : data_o = 23'b 11100111111000101111100 ;
		12'd 101 : data_o = 23'b 11100111101001110111010 ;
		12'd 102 : data_o = 23'b 11100111011010111111110 ;
		12'd 103 : data_o = 23'b 11100111001100001001000 ;
		12'd 104 : data_o = 23'b 11100110111101010010111 ;
		12'd 105 : data_o = 23'b 11100110101110011101011 ;
		12'd 106 : data_o = 23'b 11100110011111101000101 ;
		12'd 107 : data_o = 23'b 11100110010000110100100 ;
		12'd 108 : data_o = 23'b 11100110000010000001001 ;
		12'd 109 : data_o = 23'b 11100101110011001110011 ;
		12'd 110 : data_o = 23'b 11100101100100011100010 ;
		12'd 111 : data_o = 23'b 11100101010101101010111 ;
		12'd 112 : data_o = 23'b 11100101000110111010001 ;
		12'd 113 : data_o = 23'b 11100100111000001010000 ;
		12'd 114 : data_o = 23'b 11100100101001011010101 ;
		12'd 115 : data_o = 23'b 11100100011010101100000 ;
		12'd 116 : data_o = 23'b 11100100001011111101111 ;
		12'd 117 : data_o = 23'b 11100011111101010000100 ;
		12'd 118 : data_o = 23'b 11100011101110100011111 ;
		12'd 119 : data_o = 23'b 11100011011111110111111 ;
		12'd 120 : data_o = 23'b 11100011010001001100100 ;
		12'd 121 : data_o = 23'b 11100011000010100001110 ;
		12'd 122 : data_o = 23'b 11100010110011110111110 ;
		12'd 123 : data_o = 23'b 11100010100101001110011 ;
		12'd 124 : data_o = 23'b 11100010010110100101110 ;
		12'd 125 : data_o = 23'b 11100010000111111101101 ;
		12'd 126 : data_o = 23'b 11100001111001010110010 ;
		12'd 127 : data_o = 23'b 11100001101010101111101 ;
		12'd 128 : data_o = 23'b 11100001011100001001101 ;
		12'd 129 : data_o = 23'b 11100001001101100100010 ;
		12'd 130 : data_o = 23'b 11100000111110111111100 ;
		12'd 131 : data_o = 23'b 11100000110000011011100 ;
		12'd 132 : data_o = 23'b 11100000100001111000001 ;
		12'd 133 : data_o = 23'b 11100000010011010101011 ;
		12'd 134 : data_o = 23'b 11100000000100110011010 ;
		12'd 135 : data_o = 23'b 11011111110110010001111 ;
		12'd 136 : data_o = 23'b 11011111100111110001001 ;
		12'd 137 : data_o = 23'b 11011111011001010001000 ;
		12'd 138 : data_o = 23'b 11011111001010110001101 ;
		12'd 139 : data_o = 23'b 11011110111100010010111 ;
		12'd 140 : data_o = 23'b 11011110101101110100110 ;
		12'd 141 : data_o = 23'b 11011110011111010111010 ;
		12'd 142 : data_o = 23'b 11011110010000111010100 ;
		12'd 143 : data_o = 23'b 11011110000010011110010 ;
		12'd 144 : data_o = 23'b 11011101110100000010110 ;
		12'd 145 : data_o = 23'b 11011101100101101000000 ;
		12'd 146 : data_o = 23'b 11011101010111001101110 ;
		12'd 147 : data_o = 23'b 11011101001000110100010 ;
		12'd 148 : data_o = 23'b 11011100111010011011011 ;
		12'd 149 : data_o = 23'b 11011100101100000011001 ;
		12'd 150 : data_o = 23'b 11011100011101101011100 ;
		12'd 151 : data_o = 23'b 11011100001111010100101 ;
		12'd 152 : data_o = 23'b 11011100000000111110010 ;
		12'd 153 : data_o = 23'b 11011011110010101000101 ;
		12'd 154 : data_o = 23'b 11011011100100010011101 ;
		12'd 155 : data_o = 23'b 11011011010101111111010 ;
		12'd 156 : data_o = 23'b 11011011000111101011101 ;
		12'd 157 : data_o = 23'b 11011010111001011000100 ;
		12'd 158 : data_o = 23'b 11011010101011000110001 ;
		12'd 159 : data_o = 23'b 11011010011100110100011 ;
		12'd 160 : data_o = 23'b 11011010001110100011010 ;
		12'd 161 : data_o = 23'b 11011010000000010010110 ;
		12'd 162 : data_o = 23'b 11011001110010000011000 ;
		12'd 163 : data_o = 23'b 11011001100011110011110 ;
		12'd 164 : data_o = 23'b 11011001010101100101010 ;
		12'd 165 : data_o = 23'b 11011001000111010111010 ;
		12'd 166 : data_o = 23'b 11011000111001001010000 ;
		12'd 167 : data_o = 23'b 11011000101010111101011 ;
		12'd 168 : data_o = 23'b 11011000011100110001011 ;
		12'd 169 : data_o = 23'b 11011000001110100110000 ;
		12'd 170 : data_o = 23'b 11011000000000011011011 ;
		12'd 171 : data_o = 23'b 11010111110010010001010 ;
		12'd 172 : data_o = 23'b 11010111100100000111111 ;
		12'd 173 : data_o = 23'b 11010111010101111111000 ;
		12'd 174 : data_o = 23'b 11010111000111110110111 ;
		12'd 175 : data_o = 23'b 11010110111001101111011 ;
		12'd 176 : data_o = 23'b 11010110101011101000011 ;
		12'd 177 : data_o = 23'b 11010110011101100010001 ;
		12'd 178 : data_o = 23'b 11010110001111011100100 ;
		12'd 179 : data_o = 23'b 11010110000001010111100 ;
		12'd 180 : data_o = 23'b 11010101110011010011001 ;
		12'd 181 : data_o = 23'b 11010101100101001111011 ;
		12'd 182 : data_o = 23'b 11010101010111001100011 ;
		12'd 183 : data_o = 23'b 11010101001001001001111 ;
		12'd 184 : data_o = 23'b 11010100111011001000000 ;
		12'd 185 : data_o = 23'b 11010100101101000110110 ;
		12'd 186 : data_o = 23'b 11010100011111000110010 ;
		12'd 187 : data_o = 23'b 11010100010001000110010 ;
		12'd 188 : data_o = 23'b 11010100000011000110111 ;
		12'd 189 : data_o = 23'b 11010011110101001000010 ;
		12'd 190 : data_o = 23'b 11010011100111001010001 ;
		12'd 191 : data_o = 23'b 11010011011001001100110 ;
		12'd 192 : data_o = 23'b 11010011001011001111111 ;
		12'd 193 : data_o = 23'b 11010010111101010011101 ;
		12'd 194 : data_o = 23'b 11010010101111011000001 ;
		12'd 195 : data_o = 23'b 11010010100001011101001 ;
		12'd 196 : data_o = 23'b 11010010010011100010110 ;
		12'd 197 : data_o = 23'b 11010010000101101001001 ;
		12'd 198 : data_o = 23'b 11010001110111110000000 ;
		12'd 199 : data_o = 23'b 11010001101001110111100 ;
		12'd 200 : data_o = 23'b 11010001011011111111101 ;
		12'd 201 : data_o = 23'b 11010001001110001000100 ;
		12'd 202 : data_o = 23'b 11010001000000010001111 ;
		12'd 203 : data_o = 23'b 11010000110010011011111 ;
		12'd 204 : data_o = 23'b 11010000100100100110100 ;
		12'd 205 : data_o = 23'b 11010000010110110001110 ;
		12'd 206 : data_o = 23'b 11010000001000111101101 ;
		12'd 207 : data_o = 23'b 11001111111011001010000 ;
		12'd 208 : data_o = 23'b 11001111101101010111001 ;
		12'd 209 : data_o = 23'b 11001111011111100100111 ;
		12'd 210 : data_o = 23'b 11001111010001110011010 ;
		12'd 211 : data_o = 23'b 11001111000100000010001 ;
		12'd 212 : data_o = 23'b 11001110110110010001101 ;
		12'd 213 : data_o = 23'b 11001110101000100001111 ;
		12'd 214 : data_o = 23'b 11001110011010110010101 ;
		12'd 215 : data_o = 23'b 11001110001101000100000 ;
		12'd 216 : data_o = 23'b 11001101111111010110000 ;
		12'd 217 : data_o = 23'b 11001101110001101000101 ;
		12'd 218 : data_o = 23'b 11001101100011111011111 ;
		12'd 219 : data_o = 23'b 11001101010110001111101 ;
		12'd 220 : data_o = 23'b 11001101001000100100001 ;
		12'd 221 : data_o = 23'b 11001100111010111001001 ;
		12'd 222 : data_o = 23'b 11001100101101001110110 ;
		12'd 223 : data_o = 23'b 11001100011111100101001 ;
		12'd 224 : data_o = 23'b 11001100010001111100000 ;
		12'd 225 : data_o = 23'b 11001100000100010011011 ;
		12'd 226 : data_o = 23'b 11001011110110101011100 ;
		12'd 227 : data_o = 23'b 11001011101001000100001 ;
		12'd 228 : data_o = 23'b 11001011011011011101100 ;
		12'd 229 : data_o = 23'b 11001011001101110111011 ;
		12'd 230 : data_o = 23'b 11001011000000010001111 ;
		12'd 231 : data_o = 23'b 11001010110010101101000 ;
		12'd 232 : data_o = 23'b 11001010100101001000101 ;
		12'd 233 : data_o = 23'b 11001010010111100101000 ;
		12'd 234 : data_o = 23'b 11001010001010000001111 ;
		12'd 235 : data_o = 23'b 11001001111100011111011 ;
		12'd 236 : data_o = 23'b 11001001101110111101100 ;
		12'd 237 : data_o = 23'b 11001001100001011100010 ;
		12'd 238 : data_o = 23'b 11001001010011111011100 ;
		12'd 239 : data_o = 23'b 11001001000110011011011 ;
		12'd 240 : data_o = 23'b 11001000111000111011111 ;
		12'd 241 : data_o = 23'b 11001000101011011101000 ;
		12'd 242 : data_o = 23'b 11001000011101111110110 ;
		12'd 243 : data_o = 23'b 11001000010000100001000 ;
		12'd 244 : data_o = 23'b 11001000000011000011111 ;
		12'd 245 : data_o = 23'b 11000111110101100111011 ;
		12'd 246 : data_o = 23'b 11000111101000001011011 ;
		12'd 247 : data_o = 23'b 11000111011010110000001 ;
		12'd 248 : data_o = 23'b 11000111001101010101011 ;
		12'd 249 : data_o = 23'b 11000110111111111011010 ;
		12'd 250 : data_o = 23'b 11000110110010100001101 ;
		12'd 251 : data_o = 23'b 11000110100101001000110 ;
		12'd 252 : data_o = 23'b 11000110010111110000011 ;
		12'd 253 : data_o = 23'b 11000110001010011000100 ;
		12'd 254 : data_o = 23'b 11000101111101000001011 ;
		12'd 255 : data_o = 23'b 11000101101111101010110 ;
		12'd 256 : data_o = 23'b 11000101100010010100110 ;
		12'd 257 : data_o = 23'b 11000101010100111111011 ;
		12'd 258 : data_o = 23'b 11000101000111101010100 ;
		12'd 259 : data_o = 23'b 11000100111010010110010 ;
		12'd 260 : data_o = 23'b 11000100101101000010101 ;
		12'd 261 : data_o = 23'b 11000100011111101111100 ;
		12'd 262 : data_o = 23'b 11000100010010011101000 ;
		12'd 263 : data_o = 23'b 11000100000101001011001 ;
		12'd 264 : data_o = 23'b 11000011110111111001111 ;
		12'd 265 : data_o = 23'b 11000011101010101001001 ;
		12'd 266 : data_o = 23'b 11000011011101011000111 ;
		12'd 267 : data_o = 23'b 11000011010000001001011 ;
		12'd 268 : data_o = 23'b 11000011000010111010011 ;
		12'd 269 : data_o = 23'b 11000010110101101100000 ;
		12'd 270 : data_o = 23'b 11000010101000011110001 ;
		12'd 271 : data_o = 23'b 11000010011011010000111 ;
		12'd 272 : data_o = 23'b 11000010001110000100010 ;
		12'd 273 : data_o = 23'b 11000010000000111000010 ;
		12'd 274 : data_o = 23'b 11000001110011101100110 ;
		12'd 275 : data_o = 23'b 11000001100110100001110 ;
		12'd 276 : data_o = 23'b 11000001011001010111011 ;
		12'd 277 : data_o = 23'b 11000001001100001101101 ;
		12'd 278 : data_o = 23'b 11000000111111000100100 ;
		12'd 279 : data_o = 23'b 11000000110001111011111 ;
		12'd 280 : data_o = 23'b 11000000100100110011111 ;
		12'd 281 : data_o = 23'b 11000000010111101100011 ;
		12'd 282 : data_o = 23'b 11000000001010100101100 ;
		12'd 283 : data_o = 23'b 10111111111101011111001 ;
		12'd 284 : data_o = 23'b 10111111110000011001100 ;
		12'd 285 : data_o = 23'b 10111111100011010100010 ;
		12'd 286 : data_o = 23'b 10111111010110001111110 ;
		12'd 287 : data_o = 23'b 10111111001001001011101 ;
		12'd 288 : data_o = 23'b 10111110111100001000010 ;
		12'd 289 : data_o = 23'b 10111110101111000101011 ;
		12'd 290 : data_o = 23'b 10111110100010000011001 ;
		12'd 291 : data_o = 23'b 10111110010101000001011 ;
		12'd 292 : data_o = 23'b 10111110001000000000001 ;
		12'd 293 : data_o = 23'b 10111101111010111111101 ;
		12'd 294 : data_o = 23'b 10111101101101111111101 ;
		12'd 295 : data_o = 23'b 10111101100001000000001 ;
		12'd 296 : data_o = 23'b 10111101010100000001010 ;
		12'd 297 : data_o = 23'b 10111101000111000010111 ;
		12'd 298 : data_o = 23'b 10111100111010000101001 ;
		12'd 299 : data_o = 23'b 10111100101101001000000 ;
		12'd 300 : data_o = 23'b 10111100100000001011011 ;
		12'd 301 : data_o = 23'b 10111100010011001111010 ;
		12'd 302 : data_o = 23'b 10111100000110010011111 ;
		12'd 303 : data_o = 23'b 10111011111001011000111 ;
		12'd 304 : data_o = 23'b 10111011101100011110100 ;
		12'd 305 : data_o = 23'b 10111011011111100100110 ;
		12'd 306 : data_o = 23'b 10111011010010101011100 ;
		12'd 307 : data_o = 23'b 10111011000101110010111 ;
		12'd 308 : data_o = 23'b 10111010111000111010110 ;
		12'd 309 : data_o = 23'b 10111010101100000011001 ;
		12'd 310 : data_o = 23'b 10111010011111001100001 ;
		12'd 311 : data_o = 23'b 10111010010010010101110 ;
		12'd 312 : data_o = 23'b 10111010000101011111111 ;
		12'd 313 : data_o = 23'b 10111001111000101010101 ;
		12'd 314 : data_o = 23'b 10111001101011110101110 ;
		12'd 315 : data_o = 23'b 10111001011111000001101 ;
		12'd 316 : data_o = 23'b 10111001010010001110000 ;
		12'd 317 : data_o = 23'b 10111001000101011010111 ;
		12'd 318 : data_o = 23'b 10111000111000101000011 ;
		12'd 319 : data_o = 23'b 10111000101011110110011 ;
		12'd 320 : data_o = 23'b 10111000011111000101000 ;
		12'd 321 : data_o = 23'b 10111000010010010100001 ;
		12'd 322 : data_o = 23'b 10111000000101100011111 ;
		12'd 323 : data_o = 23'b 10110111111000110100001 ;
		12'd 324 : data_o = 23'b 10110111101100000100111 ;
		12'd 325 : data_o = 23'b 10110111011111010110010 ;
		12'd 326 : data_o = 23'b 10110111010010101000001 ;
		12'd 327 : data_o = 23'b 10110111000101111010101 ;
		12'd 328 : data_o = 23'b 10110110111001001101101 ;
		12'd 329 : data_o = 23'b 10110110101100100001010 ;
		12'd 330 : data_o = 23'b 10110110011111110101011 ;
		12'd 331 : data_o = 23'b 10110110010011001010000 ;
		12'd 332 : data_o = 23'b 10110110000110011111010 ;
		12'd 333 : data_o = 23'b 10110101111001110101000 ;
		12'd 334 : data_o = 23'b 10110101101101001011011 ;
		12'd 335 : data_o = 23'b 10110101100000100010001 ;
		12'd 336 : data_o = 23'b 10110101010011111001101 ;
		12'd 337 : data_o = 23'b 10110101000111010001100 ;
		12'd 338 : data_o = 23'b 10110100111010101010000 ;
		12'd 339 : data_o = 23'b 10110100101110000011001 ;
		12'd 340 : data_o = 23'b 10110100100001011100110 ;
		12'd 341 : data_o = 23'b 10110100010100110110111 ;
		12'd 342 : data_o = 23'b 10110100001000010001100 ;
		12'd 343 : data_o = 23'b 10110011111011101100110 ;
		12'd 344 : data_o = 23'b 10110011101111001000100 ;
		12'd 345 : data_o = 23'b 10110011100010100100111 ;
		12'd 346 : data_o = 23'b 10110011010110000001110 ;
		12'd 347 : data_o = 23'b 10110011001001011111001 ;
		12'd 348 : data_o = 23'b 10110010111100111101001 ;
		12'd 349 : data_o = 23'b 10110010110000011011100 ;
		12'd 350 : data_o = 23'b 10110010100011111010101 ;
		12'd 351 : data_o = 23'b 10110010010111011010001 ;
		12'd 352 : data_o = 23'b 10110010001010111010010 ;
		12'd 353 : data_o = 23'b 10110001111110011010111 ;
		12'd 354 : data_o = 23'b 10110001110001111100001 ;
		12'd 355 : data_o = 23'b 10110001100101011101110 ;
		12'd 356 : data_o = 23'b 10110001011001000000001 ;
		12'd 357 : data_o = 23'b 10110001001100100010111 ;
		12'd 358 : data_o = 23'b 10110001000000000110010 ;
		12'd 359 : data_o = 23'b 10110000110011101010001 ;
		12'd 360 : data_o = 23'b 10110000100111001110100 ;
		12'd 361 : data_o = 23'b 10110000011010110011011 ;
		12'd 362 : data_o = 23'b 10110000001110011000111 ;
		12'd 363 : data_o = 23'b 10110000000001111110111 ;
		12'd 364 : data_o = 23'b 10101111110101100101100 ;
		12'd 365 : data_o = 23'b 10101111101001001100100 ;
		12'd 366 : data_o = 23'b 10101111011100110100001 ;
		12'd 367 : data_o = 23'b 10101111010000011100010 ;
		12'd 368 : data_o = 23'b 10101111000100000101000 ;
		12'd 369 : data_o = 23'b 10101110110111101110010 ;
		12'd 370 : data_o = 23'b 10101110101011010111111 ;
		12'd 371 : data_o = 23'b 10101110011111000010010 ;
		12'd 372 : data_o = 23'b 10101110010010101101000 ;
		12'd 373 : data_o = 23'b 10101110000110011000011 ;
		12'd 374 : data_o = 23'b 10101101111010000100010 ;
		12'd 375 : data_o = 23'b 10101101101101110000101 ;
		12'd 376 : data_o = 23'b 10101101100001011101100 ;
		12'd 377 : data_o = 23'b 10101101010101001011000 ;
		12'd 378 : data_o = 23'b 10101101001000111000111 ;
		12'd 379 : data_o = 23'b 10101100111100100111011 ;
		12'd 380 : data_o = 23'b 10101100110000010110100 ;
		12'd 381 : data_o = 23'b 10101100100100000110000 ;
		12'd 382 : data_o = 23'b 10101100010111110110001 ;
		12'd 383 : data_o = 23'b 10101100001011100110101 ;
		12'd 384 : data_o = 23'b 10101011111111010111111 ;
		12'd 385 : data_o = 23'b 10101011110011001001100 ;
		12'd 386 : data_o = 23'b 10101011100110111011101 ;
		12'd 387 : data_o = 23'b 10101011011010101110011 ;
		12'd 388 : data_o = 23'b 10101011001110100001100 ;
		12'd 389 : data_o = 23'b 10101011000010010101010 ;
		12'd 390 : data_o = 23'b 10101010110110001001101 ;
		12'd 391 : data_o = 23'b 10101010101001111110011 ;
		12'd 392 : data_o = 23'b 10101010011101110011101 ;
		12'd 393 : data_o = 23'b 10101010010001101001100 ;
		12'd 394 : data_o = 23'b 10101010000101011111111 ;
		12'd 395 : data_o = 23'b 10101001111001010110110 ;
		12'd 396 : data_o = 23'b 10101001101101001110001 ;
		12'd 397 : data_o = 23'b 10101001100001000110000 ;
		12'd 398 : data_o = 23'b 10101001010100111110011 ;
		12'd 399 : data_o = 23'b 10101001001000110111011 ;
		12'd 400 : data_o = 23'b 10101000111100110000110 ;
		12'd 401 : data_o = 23'b 10101000110000101010110 ;
		12'd 402 : data_o = 23'b 10101000100100100101010 ;
		12'd 403 : data_o = 23'b 10101000011000100000010 ;
		12'd 404 : data_o = 23'b 10101000001100011011110 ;
		12'd 405 : data_o = 23'b 10101000000000010111111 ;
		12'd 406 : data_o = 23'b 10100111110100010100011 ;
		12'd 407 : data_o = 23'b 10100111101000010001100 ;
		12'd 408 : data_o = 23'b 10100111011100001111000 ;
		12'd 409 : data_o = 23'b 10100111010000001101001 ;
		12'd 410 : data_o = 23'b 10100111000100001011110 ;
		12'd 411 : data_o = 23'b 10100110111000001010111 ;
		12'd 412 : data_o = 23'b 10100110101100001010100 ;
		12'd 413 : data_o = 23'b 10100110100000001010101 ;
		12'd 414 : data_o = 23'b 10100110010100001011010 ;
		12'd 415 : data_o = 23'b 10100110001000001100011 ;
		12'd 416 : data_o = 23'b 10100101111100001110001 ;
		12'd 417 : data_o = 23'b 10100101110000010000010 ;
		12'd 418 : data_o = 23'b 10100101100100010010111 ;
		12'd 419 : data_o = 23'b 10100101011000010110001 ;
		12'd 420 : data_o = 23'b 10100101001100011001111 ;
		12'd 421 : data_o = 23'b 10100101000000011110000 ;
		12'd 422 : data_o = 23'b 10100100110100100010110 ;
		12'd 423 : data_o = 23'b 10100100101000101000000 ;
		12'd 424 : data_o = 23'b 10100100011100101101110 ;
		12'd 425 : data_o = 23'b 10100100010000110100000 ;
		12'd 426 : data_o = 23'b 10100100000100111010101 ;
		12'd 427 : data_o = 23'b 10100011111001000001111 ;
		12'd 428 : data_o = 23'b 10100011101101001001101 ;
		12'd 429 : data_o = 23'b 10100011100001010001111 ;
		12'd 430 : data_o = 23'b 10100011010101011010110 ;
		12'd 431 : data_o = 23'b 10100011001001100100000 ;
		12'd 432 : data_o = 23'b 10100010111101101101110 ;
		12'd 433 : data_o = 23'b 10100010110001111000000 ;
		12'd 434 : data_o = 23'b 10100010100110000010110 ;
		12'd 435 : data_o = 23'b 10100010011010001110000 ;
		12'd 436 : data_o = 23'b 10100010001110011001110 ;
		12'd 437 : data_o = 23'b 10100010000010100110001 ;
		12'd 438 : data_o = 23'b 10100001110110110010111 ;
		12'd 439 : data_o = 23'b 10100001101011000000001 ;
		12'd 440 : data_o = 23'b 10100001011111001101111 ;
		12'd 441 : data_o = 23'b 10100001010011011100001 ;
		12'd 442 : data_o = 23'b 10100001000111101010111 ;
		12'd 443 : data_o = 23'b 10100000111011111010001 ;
		12'd 444 : data_o = 23'b 10100000110000001001111 ;
		12'd 445 : data_o = 23'b 10100000100100011010010 ;
		12'd 446 : data_o = 23'b 10100000011000101011000 ;
		12'd 447 : data_o = 23'b 10100000001100111100010 ;
		12'd 448 : data_o = 23'b 10100000000001001110000 ;
		12'd 449 : data_o = 23'b 10011111110101100000001 ;
		12'd 450 : data_o = 23'b 10011111101001110010111 ;
		12'd 451 : data_o = 23'b 10011111011110000110001 ;
		12'd 452 : data_o = 23'b 10011111010010011001111 ;
		12'd 453 : data_o = 23'b 10011111000110101110001 ;
		12'd 454 : data_o = 23'b 10011110111011000010110 ;
		12'd 455 : data_o = 23'b 10011110101111011000000 ;
		12'd 456 : data_o = 23'b 10011110100011101101110 ;
		12'd 457 : data_o = 23'b 10011110011000000011111 ;
		12'd 458 : data_o = 23'b 10011110001100011010101 ;
		12'd 459 : data_o = 23'b 10011110000000110001110 ;
		12'd 460 : data_o = 23'b 10011101110101001001011 ;
		12'd 461 : data_o = 23'b 10011101101001100001100 ;
		12'd 462 : data_o = 23'b 10011101011101111010001 ;
		12'd 463 : data_o = 23'b 10011101010010010011010 ;
		12'd 464 : data_o = 23'b 10011101000110101100111 ;
		12'd 465 : data_o = 23'b 10011100111011000111000 ;
		12'd 466 : data_o = 23'b 10011100101111100001101 ;
		12'd 467 : data_o = 23'b 10011100100011111100110 ;
		12'd 468 : data_o = 23'b 10011100011000011000010 ;
		12'd 469 : data_o = 23'b 10011100001100110100011 ;
		12'd 470 : data_o = 23'b 10011100000001010000111 ;
		12'd 471 : data_o = 23'b 10011011110101101101111 ;
		12'd 472 : data_o = 23'b 10011011101010001011011 ;
		12'd 473 : data_o = 23'b 10011011011110101001011 ;
		12'd 474 : data_o = 23'b 10011011010011000111111 ;
		12'd 475 : data_o = 23'b 10011011000111100110111 ;
		12'd 476 : data_o = 23'b 10011010111100000110010 ;
		12'd 477 : data_o = 23'b 10011010110000100110010 ;
		12'd 478 : data_o = 23'b 10011010100101000110101 ;
		12'd 479 : data_o = 23'b 10011010011001100111100 ;
		12'd 480 : data_o = 23'b 10011010001110001000111 ;
		12'd 481 : data_o = 23'b 10011010000010101010110 ;
		12'd 482 : data_o = 23'b 10011001110111001101001 ;
		12'd 483 : data_o = 23'b 10011001101011101111111 ;
		12'd 484 : data_o = 23'b 10011001100000010011010 ;
		12'd 485 : data_o = 23'b 10011001010100110111000 ;
		12'd 486 : data_o = 23'b 10011001001001011011010 ;
		12'd 487 : data_o = 23'b 10011000111110000000000 ;
		12'd 488 : data_o = 23'b 10011000110010100101010 ;
		12'd 489 : data_o = 23'b 10011000100111001010111 ;
		12'd 490 : data_o = 23'b 10011000011011110001001 ;
		12'd 491 : data_o = 23'b 10011000010000010111110 ;
		12'd 492 : data_o = 23'b 10011000000100111110111 ;
		12'd 493 : data_o = 23'b 10010111111001100110100 ;
		12'd 494 : data_o = 23'b 10010111101110001110100 ;
		12'd 495 : data_o = 23'b 10010111100010110111001 ;
		12'd 496 : data_o = 23'b 10010111010111100000001 ;
		12'd 497 : data_o = 23'b 10010111001100001001101 ;
		12'd 498 : data_o = 23'b 10010111000000110011101 ;
		12'd 499 : data_o = 23'b 10010110110101011110001 ;
		12'd 500 : data_o = 23'b 10010110101010001001000 ;
		12'd 501 : data_o = 23'b 10010110011110110100011 ;
		12'd 502 : data_o = 23'b 10010110010011100000010 ;
		12'd 503 : data_o = 23'b 10010110001000001100101 ;
		12'd 504 : data_o = 23'b 10010101111100111001100 ;
		12'd 505 : data_o = 23'b 10010101110001100110110 ;
		12'd 506 : data_o = 23'b 10010101100110010100100 ;
		12'd 507 : data_o = 23'b 10010101011011000010110 ;
		12'd 508 : data_o = 23'b 10010101001111110001011 ;
		12'd 509 : data_o = 23'b 10010101000100100000101 ;
		12'd 510 : data_o = 23'b 10010100111001010000010 ;
		12'd 511 : data_o = 23'b 10010100101110000000011 ;
		12'd 512 : data_o = 23'b 10010100100010110000111 ;
		12'd 513 : data_o = 23'b 10010100010111100010000 ;
		12'd 514 : data_o = 23'b 10010100001100010011100 ;
		12'd 515 : data_o = 23'b 10010100000001000101100 ;
		12'd 516 : data_o = 23'b 10010011110101110111111 ;
		12'd 517 : data_o = 23'b 10010011101010101010111 ;
		12'd 518 : data_o = 23'b 10010011011111011110010 ;
		12'd 519 : data_o = 23'b 10010011010100010010000 ;
		12'd 520 : data_o = 23'b 10010011001001000110011 ;
		12'd 521 : data_o = 23'b 10010010111101111011001 ;
		12'd 522 : data_o = 23'b 10010010110010110000011 ;
		12'd 523 : data_o = 23'b 10010010100111100110001 ;
		12'd 524 : data_o = 23'b 10010010011100011100010 ;
		12'd 525 : data_o = 23'b 10010010010001010010111 ;
		12'd 526 : data_o = 23'b 10010010000110001010000 ;
		12'd 527 : data_o = 23'b 10010001111011000001100 ;
		12'd 528 : data_o = 23'b 10010001101111111001101 ;
		12'd 529 : data_o = 23'b 10010001100100110010000 ;
		12'd 530 : data_o = 23'b 10010001011001101011000 ;
		12'd 531 : data_o = 23'b 10010001001110100100011 ;
		12'd 532 : data_o = 23'b 10010001000011011110010 ;
		12'd 533 : data_o = 23'b 10010000111000011000101 ;
		12'd 534 : data_o = 23'b 10010000101101010011011 ;
		12'd 535 : data_o = 23'b 10010000100010001110101 ;
		12'd 536 : data_o = 23'b 10010000010111001010011 ;
		12'd 537 : data_o = 23'b 10010000001100000110100 ;
		12'd 538 : data_o = 23'b 10010000000001000011001 ;
		12'd 539 : data_o = 23'b 10001111110110000000010 ;
		12'd 540 : data_o = 23'b 10001111101010111101110 ;
		12'd 541 : data_o = 23'b 10001111011111111011110 ;
		12'd 542 : data_o = 23'b 10001111010100111010001 ;
		12'd 543 : data_o = 23'b 10001111001001111001001 ;
		12'd 544 : data_o = 23'b 10001110111110111000100 ;
		12'd 545 : data_o = 23'b 10001110110011111000010 ;
		12'd 546 : data_o = 23'b 10001110101000111000100 ;
		12'd 547 : data_o = 23'b 10001110011101111001010 ;
		12'd 548 : data_o = 23'b 10001110010010111010011 ;
		12'd 549 : data_o = 23'b 10001110000111111100001 ;
		12'd 550 : data_o = 23'b 10001101111100111110001 ;
		12'd 551 : data_o = 23'b 10001101110010000000110 ;
		12'd 552 : data_o = 23'b 10001101100111000011110 ;
		12'd 553 : data_o = 23'b 10001101011100000111001 ;
		12'd 554 : data_o = 23'b 10001101010001001011000 ;
		12'd 555 : data_o = 23'b 10001101000110001111011 ;
		12'd 556 : data_o = 23'b 10001100111011010100010 ;
		12'd 557 : data_o = 23'b 10001100110000011001100 ;
		12'd 558 : data_o = 23'b 10001100100101011111001 ;
		12'd 559 : data_o = 23'b 10001100011010100101010 ;
		12'd 560 : data_o = 23'b 10001100001111101011111 ;
		12'd 561 : data_o = 23'b 10001100000100110011000 ;
		12'd 562 : data_o = 23'b 10001011111001111010100 ;
		12'd 563 : data_o = 23'b 10001011101111000010011 ;
		12'd 564 : data_o = 23'b 10001011100100001010110 ;
		12'd 565 : data_o = 23'b 10001011011001010011101 ;
		12'd 566 : data_o = 23'b 10001011001110011100111 ;
		12'd 567 : data_o = 23'b 10001011000011100110101 ;
		12'd 568 : data_o = 23'b 10001010111000110000111 ;
		12'd 569 : data_o = 23'b 10001010101101111011100 ;
		12'd 570 : data_o = 23'b 10001010100011000110100 ;
		12'd 571 : data_o = 23'b 10001010011000010010001 ;
		12'd 572 : data_o = 23'b 10001010001101011110000 ;
		12'd 573 : data_o = 23'b 10001010000010101010100 ;
		12'd 574 : data_o = 23'b 10001001110111110111011 ;
		12'd 575 : data_o = 23'b 10001001101101000100101 ;
		12'd 576 : data_o = 23'b 10001001100010010010011 ;
		12'd 577 : data_o = 23'b 10001001010111100000100 ;
		12'd 578 : data_o = 23'b 10001001001100101111001 ;
		12'd 579 : data_o = 23'b 10001001000001111110010 ;
		12'd 580 : data_o = 23'b 10001000110111001101110 ;
		12'd 581 : data_o = 23'b 10001000101100011101110 ;
		12'd 582 : data_o = 23'b 10001000100001101110001 ;
		12'd 583 : data_o = 23'b 10001000010110111111000 ;
		12'd 584 : data_o = 23'b 10001000001100010000010 ;
		12'd 585 : data_o = 23'b 10001000000001100010000 ;
		12'd 586 : data_o = 23'b 10000111110110110100001 ;
		12'd 587 : data_o = 23'b 10000111101100000110110 ;
		12'd 588 : data_o = 23'b 10000111100001011001110 ;
		12'd 589 : data_o = 23'b 10000111010110101101010 ;
		12'd 590 : data_o = 23'b 10000111001100000001001 ;
		12'd 591 : data_o = 23'b 10000111000001010101100 ;
		12'd 592 : data_o = 23'b 10000110110110101010010 ;
		12'd 593 : data_o = 23'b 10000110101011111111100 ;
		12'd 594 : data_o = 23'b 10000110100001010101001 ;
		12'd 595 : data_o = 23'b 10000110010110101011010 ;
		12'd 596 : data_o = 23'b 10000110001100000001110 ;
		12'd 597 : data_o = 23'b 10000110000001011000110 ;
		12'd 598 : data_o = 23'b 10000101110110110000001 ;
		12'd 599 : data_o = 23'b 10000101101100001000000 ;
		12'd 600 : data_o = 23'b 10000101100001100000010 ;
		12'd 601 : data_o = 23'b 10000101010110111001000 ;
		12'd 602 : data_o = 23'b 10000101001100010010001 ;
		12'd 603 : data_o = 23'b 10000101000001101011101 ;
		12'd 604 : data_o = 23'b 10000100110111000101101 ;
		12'd 605 : data_o = 23'b 10000100101100100000001 ;
		12'd 606 : data_o = 23'b 10000100100001111011000 ;
		12'd 607 : data_o = 23'b 10000100010111010110010 ;
		12'd 608 : data_o = 23'b 10000100001100110010000 ;
		12'd 609 : data_o = 23'b 10000100000010001110010 ;
		12'd 610 : data_o = 23'b 10000011110111101010110 ;
		12'd 611 : data_o = 23'b 10000011101101000111111 ;
		12'd 612 : data_o = 23'b 10000011100010100101010 ;
		12'd 613 : data_o = 23'b 10000011011000000011001 ;
		12'd 614 : data_o = 23'b 10000011001101100001100 ;
		12'd 615 : data_o = 23'b 10000011000011000000010 ;
		12'd 616 : data_o = 23'b 10000010111000011111011 ;
		12'd 617 : data_o = 23'b 10000010101101111111000 ;
		12'd 618 : data_o = 23'b 10000010100011011111000 ;
		12'd 619 : data_o = 23'b 10000010011000111111100 ;
		12'd 620 : data_o = 23'b 10000010001110100000011 ;
		12'd 621 : data_o = 23'b 10000010000100000001110 ;
		12'd 622 : data_o = 23'b 10000001111001100011100 ;
		12'd 623 : data_o = 23'b 10000001101111000101101 ;
		12'd 624 : data_o = 23'b 10000001100100101000010 ;
		12'd 625 : data_o = 23'b 10000001011010001011010 ;
		12'd 626 : data_o = 23'b 10000001001111101110101 ;
		12'd 627 : data_o = 23'b 10000001000101010010100 ;
		12'd 628 : data_o = 23'b 10000000111010110110110 ;
		12'd 629 : data_o = 23'b 10000000110000011011100 ;
		12'd 630 : data_o = 23'b 10000000100110000000101 ;
		12'd 631 : data_o = 23'b 10000000011011100110010 ;
		12'd 632 : data_o = 23'b 10000000010001001100010 ;
		12'd 633 : data_o = 23'b 10000000000110110010101 ;
		12'd 634 : data_o = 23'b 01111111111100011001100 ;
		12'd 635 : data_o = 23'b 01111111110010000000110 ;
		12'd 636 : data_o = 23'b 01111111100111101000011 ;
		12'd 637 : data_o = 23'b 01111111011101010000100 ;
		12'd 638 : data_o = 23'b 01111111010010111001000 ;
		12'd 639 : data_o = 23'b 01111111001000100001111 ;
		12'd 640 : data_o = 23'b 01111110111110001011010 ;
		12'd 641 : data_o = 23'b 01111110110011110101000 ;
		12'd 642 : data_o = 23'b 01111110101001011111010 ;
		12'd 643 : data_o = 23'b 01111110011111001001111 ;
		12'd 644 : data_o = 23'b 01111110010100110100111 ;
		12'd 645 : data_o = 23'b 01111110001010100000010 ;
		12'd 646 : data_o = 23'b 01111110000000001100001 ;
		12'd 647 : data_o = 23'b 01111101110101111000100 ;
		12'd 648 : data_o = 23'b 01111101101011100101001 ;
		12'd 649 : data_o = 23'b 01111101100001010010010 ;
		12'd 650 : data_o = 23'b 01111101010110111111110 ;
		12'd 651 : data_o = 23'b 01111101001100101101110 ;
		12'd 652 : data_o = 23'b 01111101000010011100001 ;
		12'd 653 : data_o = 23'b 01111100111000001010111 ;
		12'd 654 : data_o = 23'b 01111100101101111010001 ;
		12'd 655 : data_o = 23'b 01111100100011101001110 ;
		12'd 656 : data_o = 23'b 01111100011001011001110 ;
		12'd 657 : data_o = 23'b 01111100001111001010001 ;
		12'd 658 : data_o = 23'b 01111100000100111011000 ;
		12'd 659 : data_o = 23'b 01111011111010101100010 ;
		12'd 660 : data_o = 23'b 01111011110000011110000 ;
		12'd 661 : data_o = 23'b 01111011100110010000000 ;
		12'd 662 : data_o = 23'b 01111011011100000010100 ;
		12'd 663 : data_o = 23'b 01111011010001110101100 ;
		12'd 664 : data_o = 23'b 01111011000111101000110 ;
		12'd 665 : data_o = 23'b 01111010111101011100100 ;
		12'd 666 : data_o = 23'b 01111010110011010000101 ;
		12'd 667 : data_o = 23'b 01111010101001000101010 ;
		12'd 668 : data_o = 23'b 01111010011110111010010 ;
		12'd 669 : data_o = 23'b 01111010010100101111101 ;
		12'd 670 : data_o = 23'b 01111010001010100101011 ;
		12'd 671 : data_o = 23'b 01111010000000011011101 ;
		12'd 672 : data_o = 23'b 01111001110110010010001 ;
		12'd 673 : data_o = 23'b 01111001101100001001010 ;
		12'd 674 : data_o = 23'b 01111001100010000000101 ;
		12'd 675 : data_o = 23'b 01111001010111111000100 ;
		12'd 676 : data_o = 23'b 01111001001101110000110 ;
		12'd 677 : data_o = 23'b 01111001000011101001011 ;
		12'd 678 : data_o = 23'b 01111000111001100010011 ;
		12'd 679 : data_o = 23'b 01111000101111011011111 ;
		12'd 680 : data_o = 23'b 01111000100101010101110 ;
		12'd 681 : data_o = 23'b 01111000011011010000000 ;
		12'd 682 : data_o = 23'b 01111000010001001010101 ;
		12'd 683 : data_o = 23'b 01111000000111000101110 ;
		12'd 684 : data_o = 23'b 01110111111101000001010 ;
		12'd 685 : data_o = 23'b 01110111110010111101001 ;
		12'd 686 : data_o = 23'b 01110111101000111001011 ;
		12'd 687 : data_o = 23'b 01110111011110110110001 ;
		12'd 688 : data_o = 23'b 01110111010100110011010 ;
		12'd 689 : data_o = 23'b 01110111001010110000110 ;
		12'd 690 : data_o = 23'b 01110111000000101110101 ;
		12'd 691 : data_o = 23'b 01110110110110101100111 ;
		12'd 692 : data_o = 23'b 01110110101100101011101 ;
		12'd 693 : data_o = 23'b 01110110100010101010110 ;
		12'd 694 : data_o = 23'b 01110110011000101010010 ;
		12'd 695 : data_o = 23'b 01110110001110101010010 ;
		12'd 696 : data_o = 23'b 01110110000100101010100 ;
		12'd 697 : data_o = 23'b 01110101111010101011010 ;
		12'd 698 : data_o = 23'b 01110101110000101100011 ;
		12'd 699 : data_o = 23'b 01110101100110101101111 ;
		12'd 700 : data_o = 23'b 01110101011100101111110 ;
		12'd 701 : data_o = 23'b 01110101010010110010001 ;
		12'd 702 : data_o = 23'b 01110101001000110100110 ;
		12'd 703 : data_o = 23'b 01110100111110110111111 ;
		12'd 704 : data_o = 23'b 01110100110100111011011 ;
		12'd 705 : data_o = 23'b 01110100101010111111011 ;
		12'd 706 : data_o = 23'b 01110100100001000011101 ;
		12'd 707 : data_o = 23'b 01110100010111001000011 ;
		12'd 708 : data_o = 23'b 01110100001101001101011 ;
		12'd 709 : data_o = 23'b 01110100000011010010111 ;
		12'd 710 : data_o = 23'b 01110011111001011000111 ;
		12'd 711 : data_o = 23'b 01110011101111011111001 ;
		12'd 712 : data_o = 23'b 01110011100101100101110 ;
		12'd 713 : data_o = 23'b 01110011011011101100111 ;
		12'd 714 : data_o = 23'b 01110011010001110100011 ;
		12'd 715 : data_o = 23'b 01110011000111111100010 ;
		12'd 716 : data_o = 23'b 01110010111110000100100 ;
		12'd 717 : data_o = 23'b 01110010110100001101001 ;
		12'd 718 : data_o = 23'b 01110010101010010110001 ;
		12'd 719 : data_o = 23'b 01110010100000011111101 ;
		12'd 720 : data_o = 23'b 01110010010110101001011 ;
		12'd 721 : data_o = 23'b 01110010001100110011101 ;
		12'd 722 : data_o = 23'b 01110010000010111110010 ;
		12'd 723 : data_o = 23'b 01110001111001001001010 ;
		12'd 724 : data_o = 23'b 01110001101111010100110 ;
		12'd 725 : data_o = 23'b 01110001100101100000100 ;
		12'd 726 : data_o = 23'b 01110001011011101100101 ;
		12'd 727 : data_o = 23'b 01110001010001111001010 ;
		12'd 728 : data_o = 23'b 01110001001000000110010 ;
		12'd 729 : data_o = 23'b 01110000111110010011100 ;
		12'd 730 : data_o = 23'b 01110000110100100001010 ;
		12'd 731 : data_o = 23'b 01110000101010101111011 ;
		12'd 732 : data_o = 23'b 01110000100000111110000 ;
		12'd 733 : data_o = 23'b 01110000010111001100111 ;
		12'd 734 : data_o = 23'b 01110000001101011100001 ;
		12'd 735 : data_o = 23'b 01110000000011101011111 ;
		12'd 736 : data_o = 23'b 01101111111001111011111 ;
		12'd 737 : data_o = 23'b 01101111110000001100011 ;
		12'd 738 : data_o = 23'b 01101111100110011101010 ;
		12'd 739 : data_o = 23'b 01101111011100101110100 ;
		12'd 740 : data_o = 23'b 01101111010011000000001 ;
		12'd 741 : data_o = 23'b 01101111001001010010001 ;
		12'd 742 : data_o = 23'b 01101110111111100100100 ;
		12'd 743 : data_o = 23'b 01101110110101110111010 ;
		12'd 744 : data_o = 23'b 01101110101100001010011 ;
		12'd 745 : data_o = 23'b 01101110100010011110000 ;
		12'd 746 : data_o = 23'b 01101110011000110001111 ;
		12'd 747 : data_o = 23'b 01101110001111000110010 ;
		12'd 748 : data_o = 23'b 01101110000101011010111 ;
		12'd 749 : data_o = 23'b 01101101111011110000000 ;
		12'd 750 : data_o = 23'b 01101101110010000101100 ;
		12'd 751 : data_o = 23'b 01101101101000011011010 ;
		12'd 752 : data_o = 23'b 01101101011110110001100 ;
		12'd 753 : data_o = 23'b 01101101010101001000001 ;
		12'd 754 : data_o = 23'b 01101101001011011111001 ;
		12'd 755 : data_o = 23'b 01101101000001110110100 ;
		12'd 756 : data_o = 23'b 01101100111000001110010 ;
		12'd 757 : data_o = 23'b 01101100101110100110011 ;
		12'd 758 : data_o = 23'b 01101100100100111110111 ;
		12'd 759 : data_o = 23'b 01101100011011010111111 ;
		12'd 760 : data_o = 23'b 01101100010001110001001 ;
		12'd 761 : data_o = 23'b 01101100001000001010110 ;
		12'd 762 : data_o = 23'b 01101011111110100100110 ;
		12'd 763 : data_o = 23'b 01101011110100111111010 ;
		12'd 764 : data_o = 23'b 01101011101011011010000 ;
		12'd 765 : data_o = 23'b 01101011100001110101010 ;
		12'd 766 : data_o = 23'b 01101011011000010000110 ;
		12'd 767 : data_o = 23'b 01101011001110101100101 ;
		12'd 768 : data_o = 23'b 01101011000101001001000 ;
		12'd 769 : data_o = 23'b 01101010111011100101101 ;
		12'd 770 : data_o = 23'b 01101010110010000010110 ;
		12'd 771 : data_o = 23'b 01101010101000100000001 ;
		12'd 772 : data_o = 23'b 01101010011110111110000 ;
		12'd 773 : data_o = 23'b 01101010010101011100001 ;
		12'd 774 : data_o = 23'b 01101010001011111010110 ;
		12'd 775 : data_o = 23'b 01101010000010011001101 ;
		12'd 776 : data_o = 23'b 01101001111000111001000 ;
		12'd 777 : data_o = 23'b 01101001101111011000101 ;
		12'd 778 : data_o = 23'b 01101001100101111000110 ;
		12'd 779 : data_o = 23'b 01101001011100011001010 ;
		12'd 780 : data_o = 23'b 01101001010010111010000 ;
		12'd 781 : data_o = 23'b 01101001001001011011010 ;
		12'd 782 : data_o = 23'b 01101000111111111100110 ;
		12'd 783 : data_o = 23'b 01101000110110011110101 ;
		12'd 784 : data_o = 23'b 01101000101101000001000 ;
		12'd 785 : data_o = 23'b 01101000100011100011101 ;
		12'd 786 : data_o = 23'b 01101000011010000110110 ;
		12'd 787 : data_o = 23'b 01101000010000101010001 ;
		12'd 788 : data_o = 23'b 01101000000111001101111 ;
		12'd 789 : data_o = 23'b 01100111111101110010001 ;
		12'd 790 : data_o = 23'b 01100111110100010110101 ;
		12'd 791 : data_o = 23'b 01100111101010111011100 ;
		12'd 792 : data_o = 23'b 01100111100001100000110 ;
		12'd 793 : data_o = 23'b 01100111011000000110100 ;
		12'd 794 : data_o = 23'b 01100111001110101100100 ;
		12'd 795 : data_o = 23'b 01100111000101010010111 ;
		12'd 796 : data_o = 23'b 01100110111011111001101 ;
		12'd 797 : data_o = 23'b 01100110110010100000110 ;
		12'd 798 : data_o = 23'b 01100110101001001000010 ;
		12'd 799 : data_o = 23'b 01100110011111110000000 ;
		12'd 800 : data_o = 23'b 01100110010110011000010 ;
		12'd 801 : data_o = 23'b 01100110001101000000111 ;
		12'd 802 : data_o = 23'b 01100110000011101001111 ;
		12'd 803 : data_o = 23'b 01100101111010010011001 ;
		12'd 804 : data_o = 23'b 01100101110000111100111 ;
		12'd 805 : data_o = 23'b 01100101100111100110111 ;
		12'd 806 : data_o = 23'b 01100101011110010001011 ;
		12'd 807 : data_o = 23'b 01100101010100111100001 ;
		12'd 808 : data_o = 23'b 01100101001011100111010 ;
		12'd 809 : data_o = 23'b 01100101000010010010110 ;
		12'd 810 : data_o = 23'b 01100100111000111110110 ;
		12'd 811 : data_o = 23'b 01100100101111101011000 ;
		12'd 812 : data_o = 23'b 01100100100110010111100 ;
		12'd 813 : data_o = 23'b 01100100011101000100100 ;
		12'd 814 : data_o = 23'b 01100100010011110001111 ;
		12'd 815 : data_o = 23'b 01100100001010011111101 ;
		12'd 816 : data_o = 23'b 01100100000001001101101 ;
		12'd 817 : data_o = 23'b 01100011110111111100001 ;
		12'd 818 : data_o = 23'b 01100011101110101010111 ;
		12'd 819 : data_o = 23'b 01100011100101011010000 ;
		12'd 820 : data_o = 23'b 01100011011100001001100 ;
		12'd 821 : data_o = 23'b 01100011010010111001011 ;
		12'd 822 : data_o = 23'b 01100011001001101001101 ;
		12'd 823 : data_o = 23'b 01100011000000011010010 ;
		12'd 824 : data_o = 23'b 01100010110111001011010 ;
		12'd 825 : data_o = 23'b 01100010101101111100100 ;
		12'd 826 : data_o = 23'b 01100010100100101110010 ;
		12'd 827 : data_o = 23'b 01100010011011100000010 ;
		12'd 828 : data_o = 23'b 01100010010010010010101 ;
		12'd 829 : data_o = 23'b 01100010001001000101011 ;
		12'd 830 : data_o = 23'b 01100001111111111000100 ;
		12'd 831 : data_o = 23'b 01100001110110101100000 ;
		12'd 832 : data_o = 23'b 01100001101101011111111 ;
		12'd 833 : data_o = 23'b 01100001100100010100000 ;
		12'd 834 : data_o = 23'b 01100001011011001000101 ;
		12'd 835 : data_o = 23'b 01100001010001111101100 ;
		12'd 836 : data_o = 23'b 01100001001000110010110 ;
		12'd 837 : data_o = 23'b 01100000111111101000011 ;
		12'd 838 : data_o = 23'b 01100000110110011110011 ;
		12'd 839 : data_o = 23'b 01100000101101010100101 ;
		12'd 840 : data_o = 23'b 01100000100100001011011 ;
		12'd 841 : data_o = 23'b 01100000011011000010011 ;
		12'd 842 : data_o = 23'b 01100000010001111001111 ;
		12'd 843 : data_o = 23'b 01100000001000110001101 ;
		12'd 844 : data_o = 23'b 01011111111111101001101 ;
		12'd 845 : data_o = 23'b 01011111110110100010001 ;
		12'd 846 : data_o = 23'b 01011111101101011011000 ;
		12'd 847 : data_o = 23'b 01011111100100010100001 ;
		12'd 848 : data_o = 23'b 01011111011011001101101 ;
		12'd 849 : data_o = 23'b 01011111010010000111100 ;
		12'd 850 : data_o = 23'b 01011111001001000001110 ;
		12'd 851 : data_o = 23'b 01011110111111111100011 ;
		12'd 852 : data_o = 23'b 01011110110110110111010 ;
		12'd 853 : data_o = 23'b 01011110101101110010101 ;
		12'd 854 : data_o = 23'b 01011110100100101110010 ;
		12'd 855 : data_o = 23'b 01011110011011101010010 ;
		12'd 856 : data_o = 23'b 01011110010010100110101 ;
		12'd 857 : data_o = 23'b 01011110001001100011010 ;
		12'd 858 : data_o = 23'b 01011110000000100000011 ;
		12'd 859 : data_o = 23'b 01011101110111011101110 ;
		12'd 860 : data_o = 23'b 01011101101110011011100 ;
		12'd 861 : data_o = 23'b 01011101100101011001100 ;
		12'd 862 : data_o = 23'b 01011101011100011000000 ;
		12'd 863 : data_o = 23'b 01011101010011010110110 ;
		12'd 864 : data_o = 23'b 01011101001010010110000 ;
		12'd 865 : data_o = 23'b 01011101000001010101100 ;
		12'd 866 : data_o = 23'b 01011100111000010101010 ;
		12'd 867 : data_o = 23'b 01011100101111010101100 ;
		12'd 868 : data_o = 23'b 01011100100110010110000 ;
		12'd 869 : data_o = 23'b 01011100011101010110111 ;
		12'd 870 : data_o = 23'b 01011100010100011000001 ;
		12'd 871 : data_o = 23'b 01011100001011011001110 ;
		12'd 872 : data_o = 23'b 01011100000010011011101 ;
		12'd 873 : data_o = 23'b 01011011111001011101111 ;
		12'd 874 : data_o = 23'b 01011011110000100000100 ;
		12'd 875 : data_o = 23'b 01011011100111100011100 ;
		12'd 876 : data_o = 23'b 01011011011110100110111 ;
		12'd 877 : data_o = 23'b 01011011010101101010100 ;
		12'd 878 : data_o = 23'b 01011011001100101110100 ;
		12'd 879 : data_o = 23'b 01011011000011110010111 ;
		12'd 880 : data_o = 23'b 01011010111010110111100 ;
		12'd 881 : data_o = 23'b 01011010110001111100100 ;
		12'd 882 : data_o = 23'b 01011010101001000010000 ;
		12'd 883 : data_o = 23'b 01011010100000000111101 ;
		12'd 884 : data_o = 23'b 01011010010111001101110 ;
		12'd 885 : data_o = 23'b 01011010001110010100001 ;
		12'd 886 : data_o = 23'b 01011010000101011010111 ;
		12'd 887 : data_o = 23'b 01011001111100100010000 ;
		12'd 888 : data_o = 23'b 01011001110011101001100 ;
		12'd 889 : data_o = 23'b 01011001101010110001010 ;
		12'd 890 : data_o = 23'b 01011001100001111001011 ;
		12'd 891 : data_o = 23'b 01011001011001000001110 ;
		12'd 892 : data_o = 23'b 01011001010000001010101 ;
		12'd 893 : data_o = 23'b 01011001000111010011110 ;
		12'd 894 : data_o = 23'b 01011000111110011101010 ;
		12'd 895 : data_o = 23'b 01011000110101100111001 ;
		12'd 896 : data_o = 23'b 01011000101100110001010 ;
		12'd 897 : data_o = 23'b 01011000100011111011110 ;
		12'd 898 : data_o = 23'b 01011000011011000110101 ;
		12'd 899 : data_o = 23'b 01011000010010010001110 ;
		12'd 900 : data_o = 23'b 01011000001001011101011 ;
		12'd 901 : data_o = 23'b 01011000000000101001010 ;
		12'd 902 : data_o = 23'b 01010111110111110101011 ;
		12'd 903 : data_o = 23'b 01010111101111000010000 ;
		12'd 904 : data_o = 23'b 01010111100110001110111 ;
		12'd 905 : data_o = 23'b 01010111011101011100000 ;
		12'd 906 : data_o = 23'b 01010111010100101001101 ;
		12'd 907 : data_o = 23'b 01010111001011110111100 ;
		12'd 908 : data_o = 23'b 01010111000011000101110 ;
		12'd 909 : data_o = 23'b 01010110111010010100010 ;
		12'd 910 : data_o = 23'b 01010110110001100011010 ;
		12'd 911 : data_o = 23'b 01010110101000110010011 ;
		12'd 912 : data_o = 23'b 01010110100000000010000 ;
		12'd 913 : data_o = 23'b 01010110010111010001111 ;
		12'd 914 : data_o = 23'b 01010110001110100010001 ;
		12'd 915 : data_o = 23'b 01010110000101110010110 ;
		12'd 916 : data_o = 23'b 01010101111101000011101 ;
		12'd 917 : data_o = 23'b 01010101110100010100111 ;
		12'd 918 : data_o = 23'b 01010101101011100110100 ;
		12'd 919 : data_o = 23'b 01010101100010111000011 ;
		12'd 920 : data_o = 23'b 01010101011010001010101 ;
		12'd 921 : data_o = 23'b 01010101010001011101010 ;
		12'd 922 : data_o = 23'b 01010101001000110000001 ;
		12'd 923 : data_o = 23'b 01010101000000000011011 ;
		12'd 924 : data_o = 23'b 01010100110111010111000 ;
		12'd 925 : data_o = 23'b 01010100101110101010111 ;
		12'd 926 : data_o = 23'b 01010100100101111111001 ;
		12'd 927 : data_o = 23'b 01010100011101010011110 ;
		12'd 928 : data_o = 23'b 01010100010100101000101 ;
		12'd 929 : data_o = 23'b 01010100001011111101111 ;
		12'd 930 : data_o = 23'b 01010100000011010011100 ;
		12'd 931 : data_o = 23'b 01010011111010101001011 ;
		12'd 932 : data_o = 23'b 01010011110001111111101 ;
		12'd 933 : data_o = 23'b 01010011101001010110010 ;
		12'd 934 : data_o = 23'b 01010011100000101101001 ;
		12'd 935 : data_o = 23'b 01010011011000000100011 ;
		12'd 936 : data_o = 23'b 01010011001111011011111 ;
		12'd 937 : data_o = 23'b 01010011000110110011110 ;
		12'd 938 : data_o = 23'b 01010010111110001100000 ;
		12'd 939 : data_o = 23'b 01010010110101100100100 ;
		12'd 940 : data_o = 23'b 01010010101100111101011 ;
		12'd 941 : data_o = 23'b 01010010100100010110101 ;
		12'd 942 : data_o = 23'b 01010010011011110000001 ;
		12'd 943 : data_o = 23'b 01010010010011001010000 ;
		12'd 944 : data_o = 23'b 01010010001010100100001 ;
		12'd 945 : data_o = 23'b 01010010000001111110110 ;
		12'd 946 : data_o = 23'b 01010001111001011001100 ;
		12'd 947 : data_o = 23'b 01010001110000110100110 ;
		12'd 948 : data_o = 23'b 01010001101000010000010 ;
		12'd 949 : data_o = 23'b 01010001011111101100000 ;
		12'd 950 : data_o = 23'b 01010001010111001000001 ;
		12'd 951 : data_o = 23'b 01010001001110100100101 ;
		12'd 952 : data_o = 23'b 01010001000110000001011 ;
		12'd 953 : data_o = 23'b 01010000111101011110100 ;
		12'd 954 : data_o = 23'b 01010000110100111100000 ;
		12'd 955 : data_o = 23'b 01010000101100011001110 ;
		12'd 956 : data_o = 23'b 01010000100011110111111 ;
		12'd 957 : data_o = 23'b 01010000011011010110010 ;
		12'd 958 : data_o = 23'b 01010000010010110101000 ;
		12'd 959 : data_o = 23'b 01010000001010010100000 ;
		12'd 960 : data_o = 23'b 01010000000001110011100 ;
		12'd 961 : data_o = 23'b 01001111111001010011001 ;
		12'd 962 : data_o = 23'b 01001111110000110011010 ;
		12'd 963 : data_o = 23'b 01001111101000010011100 ;
		12'd 964 : data_o = 23'b 01001111011111110100010 ;
		12'd 965 : data_o = 23'b 01001111010111010101010 ;
		12'd 966 : data_o = 23'b 01001111001110110110100 ;
		12'd 967 : data_o = 23'b 01001111000110011000010 ;
		12'd 968 : data_o = 23'b 01001110111101111010001 ;
		12'd 969 : data_o = 23'b 01001110110101011100100 ;
		12'd 970 : data_o = 23'b 01001110101100111111000 ;
		12'd 971 : data_o = 23'b 01001110100100100010000 ;
		12'd 972 : data_o = 23'b 01001110011100000101010 ;
		12'd 973 : data_o = 23'b 01001110010011101000110 ;
		12'd 974 : data_o = 23'b 01001110001011001100101 ;
		12'd 975 : data_o = 23'b 01001110000010110000111 ;
		12'd 976 : data_o = 23'b 01001101111010010101011 ;
		12'd 977 : data_o = 23'b 01001101110001111010010 ;
		12'd 978 : data_o = 23'b 01001101101001011111011 ;
		12'd 979 : data_o = 23'b 01001101100001000100111 ;
		12'd 980 : data_o = 23'b 01001101011000101010110 ;
		12'd 981 : data_o = 23'b 01001101010000010000111 ;
		12'd 982 : data_o = 23'b 01001101000111110111010 ;
		12'd 983 : data_o = 23'b 01001100111111011110000 ;
		12'd 984 : data_o = 23'b 01001100110111000101001 ;
		12'd 985 : data_o = 23'b 01001100101110101100100 ;
		12'd 986 : data_o = 23'b 01001100100110010100001 ;
		12'd 987 : data_o = 23'b 01001100011101111100010 ;
		12'd 988 : data_o = 23'b 01001100010101100100100 ;
		12'd 989 : data_o = 23'b 01001100001101001101001 ;
		12'd 990 : data_o = 23'b 01001100000100110110001 ;
		12'd 991 : data_o = 23'b 01001011111100011111100 ;
		12'd 992 : data_o = 23'b 01001011110100001001000 ;
		12'd 993 : data_o = 23'b 01001011101011110011000 ;
		12'd 994 : data_o = 23'b 01001011100011011101001 ;
		12'd 995 : data_o = 23'b 01001011011011000111110 ;
		12'd 996 : data_o = 23'b 01001011010010110010101 ;
		12'd 997 : data_o = 23'b 01001011001010011101110 ;
		12'd 998 : data_o = 23'b 01001011000010001001010 ;
		12'd 999 : data_o = 23'b 01001010111001110101000 ;
		12'd 1000 : data_o = 23'b 01001010110001100001001 ;
		12'd 1001 : data_o = 23'b 01001010101001001101101 ;
		12'd 1002 : data_o = 23'b 01001010100000111010011 ;
		12'd 1003 : data_o = 23'b 01001010011000100111011 ;
		12'd 1004 : data_o = 23'b 01001010010000010100110 ;
		12'd 1005 : data_o = 23'b 01001010001000000010011 ;
		12'd 1006 : data_o = 23'b 01001001111111110000011 ;
		12'd 1007 : data_o = 23'b 01001001110111011110110 ;
		12'd 1008 : data_o = 23'b 01001001101111001101010 ;
		12'd 1009 : data_o = 23'b 01001001100110111100010 ;
		12'd 1010 : data_o = 23'b 01001001011110101011100 ;
		12'd 1011 : data_o = 23'b 01001001010110011011000 ;
		12'd 1012 : data_o = 23'b 01001001001110001010111 ;
		12'd 1013 : data_o = 23'b 01001001000101111011000 ;
		12'd 1014 : data_o = 23'b 01001000111101101011100 ;
		12'd 1015 : data_o = 23'b 01001000110101011100010 ;
		12'd 1016 : data_o = 23'b 01001000101101001101011 ;
		12'd 1017 : data_o = 23'b 01001000100100111110110 ;
		12'd 1018 : data_o = 23'b 01001000011100110000100 ;
		12'd 1019 : data_o = 23'b 01001000010100100010100 ;
		12'd 1020 : data_o = 23'b 01001000001100010100111 ;
		12'd 1021 : data_o = 23'b 01001000000100000111100 ;
		12'd 1022 : data_o = 23'b 01000111111011111010011 ;
		12'd 1023 : data_o = 23'b 01000111110011101101101 ;
		12'd 1024 : data_o = 23'b 01000111101011100001010 ;
		12'd 1025 : data_o = 23'b 01000111100011010101001 ;
		12'd 1026 : data_o = 23'b 01000111011011001001010 ;
		12'd 1027 : data_o = 23'b 01000111010010111101110 ;
		12'd 1028 : data_o = 23'b 01000111001010110010100 ;
		12'd 1029 : data_o = 23'b 01000111000010100111101 ;
		12'd 1030 : data_o = 23'b 01000110111010011101000 ;
		12'd 1031 : data_o = 23'b 01000110110010010010110 ;
		12'd 1032 : data_o = 23'b 01000110101010001000110 ;
		12'd 1033 : data_o = 23'b 01000110100001111111000 ;
		12'd 1034 : data_o = 23'b 01000110011001110101101 ;
		12'd 1035 : data_o = 23'b 01000110010001101100101 ;
		12'd 1036 : data_o = 23'b 01000110001001100011110 ;
		12'd 1037 : data_o = 23'b 01000110000001011011011 ;
		12'd 1038 : data_o = 23'b 01000101111001010011001 ;
		12'd 1039 : data_o = 23'b 01000101110001001011011 ;
		12'd 1040 : data_o = 23'b 01000101101001000011110 ;
		12'd 1041 : data_o = 23'b 01000101100000111100100 ;
		12'd 1042 : data_o = 23'b 01000101011000110101101 ;
		12'd 1043 : data_o = 23'b 01000101010000101110111 ;
		12'd 1044 : data_o = 23'b 01000101001000101000101 ;
		12'd 1045 : data_o = 23'b 01000101000000100010100 ;
		12'd 1046 : data_o = 23'b 01000100111000011100110 ;
		12'd 1047 : data_o = 23'b 01000100110000010111011 ;
		12'd 1048 : data_o = 23'b 01000100101000010010010 ;
		12'd 1049 : data_o = 23'b 01000100100000001101011 ;
		12'd 1050 : data_o = 23'b 01000100011000001000111 ;
		12'd 1051 : data_o = 23'b 01000100010000000100101 ;
		12'd 1052 : data_o = 23'b 01000100001000000000110 ;
		12'd 1053 : data_o = 23'b 01000011111111111101001 ;
		12'd 1054 : data_o = 23'b 01000011110111111001110 ;
		12'd 1055 : data_o = 23'b 01000011101111110110110 ;
		12'd 1056 : data_o = 23'b 01000011100111110100000 ;
		12'd 1057 : data_o = 23'b 01000011011111110001100 ;
		12'd 1058 : data_o = 23'b 01000011010111101111011 ;
		12'd 1059 : data_o = 23'b 01000011001111101101101 ;
		12'd 1060 : data_o = 23'b 01000011000111101100001 ;
		12'd 1061 : data_o = 23'b 01000010111111101010111 ;
		12'd 1062 : data_o = 23'b 01000010110111101001111 ;
		12'd 1063 : data_o = 23'b 01000010101111101001010 ;
		12'd 1064 : data_o = 23'b 01000010100111101000111 ;
		12'd 1065 : data_o = 23'b 01000010011111101000111 ;
		12'd 1066 : data_o = 23'b 01000010010111101001001 ;
		12'd 1067 : data_o = 23'b 01000010001111101001110 ;
		12'd 1068 : data_o = 23'b 01000010000111101010100 ;
		12'd 1069 : data_o = 23'b 01000001111111101011110 ;
		12'd 1070 : data_o = 23'b 01000001110111101101001 ;
		12'd 1071 : data_o = 23'b 01000001101111101110111 ;
		12'd 1072 : data_o = 23'b 01000001100111110000111 ;
		12'd 1073 : data_o = 23'b 01000001011111110011010 ;
		12'd 1074 : data_o = 23'b 01000001010111110101111 ;
		12'd 1075 : data_o = 23'b 01000001001111111000110 ;
		12'd 1076 : data_o = 23'b 01000001000111111100000 ;
		12'd 1077 : data_o = 23'b 01000000111111111111100 ;
		12'd 1078 : data_o = 23'b 01000000111000000011011 ;
		12'd 1079 : data_o = 23'b 01000000110000000111100 ;
		12'd 1080 : data_o = 23'b 01000000101000001011111 ;
		12'd 1081 : data_o = 23'b 01000000100000010000100 ;
		12'd 1082 : data_o = 23'b 01000000011000010101100 ;
		12'd 1083 : data_o = 23'b 01000000010000011010110 ;
		12'd 1084 : data_o = 23'b 01000000001000100000011 ;
		12'd 1085 : data_o = 23'b 01000000000000100110010 ;
		12'd 1086 : data_o = 23'b 00111111111000101100011 ;
		12'd 1087 : data_o = 23'b 00111111110000110010111 ;
		12'd 1088 : data_o = 23'b 00111111101000111001101 ;
		12'd 1089 : data_o = 23'b 00111111100001000000101 ;
		12'd 1090 : data_o = 23'b 00111111011001001000000 ;
		12'd 1091 : data_o = 23'b 00111111010001001111101 ;
		12'd 1092 : data_o = 23'b 00111111001001010111100 ;
		12'd 1093 : data_o = 23'b 00111111000001011111110 ;
		12'd 1094 : data_o = 23'b 00111110111001101000010 ;
		12'd 1095 : data_o = 23'b 00111110110001110001000 ;
		12'd 1096 : data_o = 23'b 00111110101001111010001 ;
		12'd 1097 : data_o = 23'b 00111110100010000011100 ;
		12'd 1098 : data_o = 23'b 00111110011010001101001 ;
		12'd 1099 : data_o = 23'b 00111110010010010111000 ;
		12'd 1100 : data_o = 23'b 00111110001010100001010 ;
		12'd 1101 : data_o = 23'b 00111110000010101011110 ;
		12'd 1102 : data_o = 23'b 00111101111010110110101 ;
		12'd 1103 : data_o = 23'b 00111101110011000001110 ;
		12'd 1104 : data_o = 23'b 00111101101011001101001 ;
		12'd 1105 : data_o = 23'b 00111101100011011000111 ;
		12'd 1106 : data_o = 23'b 00111101011011100100110 ;
		12'd 1107 : data_o = 23'b 00111101010011110001000 ;
		12'd 1108 : data_o = 23'b 00111101001011111101101 ;
		12'd 1109 : data_o = 23'b 00111101000100001010011 ;
		12'd 1110 : data_o = 23'b 00111100111100010111100 ;
		12'd 1111 : data_o = 23'b 00111100110100100101000 ;
		12'd 1112 : data_o = 23'b 00111100101100110010101 ;
		12'd 1113 : data_o = 23'b 00111100100101000000101 ;
		12'd 1114 : data_o = 23'b 00111100011101001110111 ;
		12'd 1115 : data_o = 23'b 00111100010101011101100 ;
		12'd 1116 : data_o = 23'b 00111100001101101100011 ;
		12'd 1117 : data_o = 23'b 00111100000101111011100 ;
		12'd 1118 : data_o = 23'b 00111011111110001010111 ;
		12'd 1119 : data_o = 23'b 00111011110110011010101 ;
		12'd 1120 : data_o = 23'b 00111011101110101010101 ;
		12'd 1121 : data_o = 23'b 00111011100110111010111 ;
		12'd 1122 : data_o = 23'b 00111011011111001011011 ;
		12'd 1123 : data_o = 23'b 00111011010111011100010 ;
		12'd 1124 : data_o = 23'b 00111011001111101101011 ;
		12'd 1125 : data_o = 23'b 00111011000111111110110 ;
		12'd 1126 : data_o = 23'b 00111011000000010000100 ;
		12'd 1127 : data_o = 23'b 00111010111000100010100 ;
		12'd 1128 : data_o = 23'b 00111010110000110100110 ;
		12'd 1129 : data_o = 23'b 00111010101001000111010 ;
		12'd 1130 : data_o = 23'b 00111010100001011010001 ;
		12'd 1131 : data_o = 23'b 00111010011001101101010 ;
		12'd 1132 : data_o = 23'b 00111010010010000000101 ;
		12'd 1133 : data_o = 23'b 00111010001010010100010 ;
		12'd 1134 : data_o = 23'b 00111010000010101000010 ;
		12'd 1135 : data_o = 23'b 00111001111010111100100 ;
		12'd 1136 : data_o = 23'b 00111001110011010001000 ;
		12'd 1137 : data_o = 23'b 00111001101011100101111 ;
		12'd 1138 : data_o = 23'b 00111001100011111010111 ;
		12'd 1139 : data_o = 23'b 00111001011100010000010 ;
		12'd 1140 : data_o = 23'b 00111001010100100101111 ;
		12'd 1141 : data_o = 23'b 00111001001100111011111 ;
		12'd 1142 : data_o = 23'b 00111001000101010010001 ;
		12'd 1143 : data_o = 23'b 00111000111101101000101 ;
		12'd 1144 : data_o = 23'b 00111000110101111111011 ;
		12'd 1145 : data_o = 23'b 00111000101110010110011 ;
		12'd 1146 : data_o = 23'b 00111000100110101101110 ;
		12'd 1147 : data_o = 23'b 00111000011111000101011 ;
		12'd 1148 : data_o = 23'b 00111000010111011101010 ;
		12'd 1149 : data_o = 23'b 00111000001111110101011 ;
		12'd 1150 : data_o = 23'b 00111000001000001101111 ;
		12'd 1151 : data_o = 23'b 00111000000000100110101 ;
		12'd 1152 : data_o = 23'b 00110111111000111111101 ;
		12'd 1153 : data_o = 23'b 00110111110001011000111 ;
		12'd 1154 : data_o = 23'b 00110111101001110010100 ;
		12'd 1155 : data_o = 23'b 00110111100010001100010 ;
		12'd 1156 : data_o = 23'b 00110111011010100110011 ;
		12'd 1157 : data_o = 23'b 00110111010011000000110 ;
		12'd 1158 : data_o = 23'b 00110111001011011011100 ;
		12'd 1159 : data_o = 23'b 00110111000011110110011 ;
		12'd 1160 : data_o = 23'b 00110110111100010001101 ;
		12'd 1161 : data_o = 23'b 00110110110100101101001 ;
		12'd 1162 : data_o = 23'b 00110110101101001001000 ;
		12'd 1163 : data_o = 23'b 00110110100101100101000 ;
		12'd 1164 : data_o = 23'b 00110110011110000001011 ;
		12'd 1165 : data_o = 23'b 00110110010110011110000 ;
		12'd 1166 : data_o = 23'b 00110110001110111010111 ;
		12'd 1167 : data_o = 23'b 00110110000111011000000 ;
		12'd 1168 : data_o = 23'b 00110101111111110101011 ;
		12'd 1169 : data_o = 23'b 00110101111000010011001 ;
		12'd 1170 : data_o = 23'b 00110101110000110001001 ;
		12'd 1171 : data_o = 23'b 00110101101001001111011 ;
		12'd 1172 : data_o = 23'b 00110101100001101101111 ;
		12'd 1173 : data_o = 23'b 00110101011010001100110 ;
		12'd 1174 : data_o = 23'b 00110101010010101011110 ;
		12'd 1175 : data_o = 23'b 00110101001011001011001 ;
		12'd 1176 : data_o = 23'b 00110101000011101010110 ;
		12'd 1177 : data_o = 23'b 00110100111100001010101 ;
		12'd 1178 : data_o = 23'b 00110100110100101010111 ;
		12'd 1179 : data_o = 23'b 00110100101101001011010 ;
		12'd 1180 : data_o = 23'b 00110100100101101100000 ;
		12'd 1181 : data_o = 23'b 00110100011110001101000 ;
		12'd 1182 : data_o = 23'b 00110100010110101110010 ;
		12'd 1183 : data_o = 23'b 00110100001111001111111 ;
		12'd 1184 : data_o = 23'b 00110100000111110001101 ;
		12'd 1185 : data_o = 23'b 00110100000000010011110 ;
		12'd 1186 : data_o = 23'b 00110011111000110110000 ;
		12'd 1187 : data_o = 23'b 00110011110001011000101 ;
		12'd 1188 : data_o = 23'b 00110011101001111011101 ;
		12'd 1189 : data_o = 23'b 00110011100010011110110 ;
		12'd 1190 : data_o = 23'b 00110011011011000010001 ;
		12'd 1191 : data_o = 23'b 00110011010011100101111 ;
		12'd 1192 : data_o = 23'b 00110011001100001001111 ;
		12'd 1193 : data_o = 23'b 00110011000100101110001 ;
		12'd 1194 : data_o = 23'b 00110010111101010010101 ;
		12'd 1195 : data_o = 23'b 00110010110101110111011 ;
		12'd 1196 : data_o = 23'b 00110010101110011100100 ;
		12'd 1197 : data_o = 23'b 00110010100111000001110 ;
		12'd 1198 : data_o = 23'b 00110010011111100111011 ;
		12'd 1199 : data_o = 23'b 00110010011000001101010 ;
		12'd 1200 : data_o = 23'b 00110010010000110011011 ;
		12'd 1201 : data_o = 23'b 00110010001001011001110 ;
		12'd 1202 : data_o = 23'b 00110010000010000000011 ;
		12'd 1203 : data_o = 23'b 00110001111010100111011 ;
		12'd 1204 : data_o = 23'b 00110001110011001110101 ;
		12'd 1205 : data_o = 23'b 00110001101011110110000 ;
		12'd 1206 : data_o = 23'b 00110001100100011101110 ;
		12'd 1207 : data_o = 23'b 00110001011101000101110 ;
		12'd 1208 : data_o = 23'b 00110001010101101110000 ;
		12'd 1209 : data_o = 23'b 00110001001110010110101 ;
		12'd 1210 : data_o = 23'b 00110001000110111111011 ;
		12'd 1211 : data_o = 23'b 00110000111111101000100 ;
		12'd 1212 : data_o = 23'b 00110000111000010001110 ;
		12'd 1213 : data_o = 23'b 00110000110000111011011 ;
		12'd 1214 : data_o = 23'b 00110000101001100101010 ;
		12'd 1215 : data_o = 23'b 00110000100010001111011 ;
		12'd 1216 : data_o = 23'b 00110000011010111001111 ;
		12'd 1217 : data_o = 23'b 00110000010011100100100 ;
		12'd 1218 : data_o = 23'b 00110000001100001111011 ;
		12'd 1219 : data_o = 23'b 00110000000100111010101 ;
		12'd 1220 : data_o = 23'b 00101111111101100110001 ;
		12'd 1221 : data_o = 23'b 00101111110110010001110 ;
		12'd 1222 : data_o = 23'b 00101111101110111101110 ;
		12'd 1223 : data_o = 23'b 00101111100111101010000 ;
		12'd 1224 : data_o = 23'b 00101111100000010110100 ;
		12'd 1225 : data_o = 23'b 00101111011001000011011 ;
		12'd 1226 : data_o = 23'b 00101111010001110000011 ;
		12'd 1227 : data_o = 23'b 00101111001010011101101 ;
		12'd 1228 : data_o = 23'b 00101111000011001011010 ;
		12'd 1229 : data_o = 23'b 00101110111011111001001 ;
		12'd 1230 : data_o = 23'b 00101110110100100111001 ;
		12'd 1231 : data_o = 23'b 00101110101101010101100 ;
		12'd 1232 : data_o = 23'b 00101110100110000100001 ;
		12'd 1233 : data_o = 23'b 00101110011110110011000 ;
		12'd 1234 : data_o = 23'b 00101110010111100010001 ;
		12'd 1235 : data_o = 23'b 00101110010000010001100 ;
		12'd 1236 : data_o = 23'b 00101110001001000001010 ;
		12'd 1237 : data_o = 23'b 00101110000001110001001 ;
		12'd 1238 : data_o = 23'b 00101101111010100001011 ;
		12'd 1239 : data_o = 23'b 00101101110011010001110 ;
		12'd 1240 : data_o = 23'b 00101101101100000010100 ;
		12'd 1241 : data_o = 23'b 00101101100100110011100 ;
		12'd 1242 : data_o = 23'b 00101101011101100100110 ;
		12'd 1243 : data_o = 23'b 00101101010110010110001 ;
		12'd 1244 : data_o = 23'b 00101101001111000111111 ;
		12'd 1245 : data_o = 23'b 00101101000111111010000 ;
		12'd 1246 : data_o = 23'b 00101101000000101100010 ;
		12'd 1247 : data_o = 23'b 00101100111001011110110 ;
		12'd 1248 : data_o = 23'b 00101100110010010001100 ;
		12'd 1249 : data_o = 23'b 00101100101011000100101 ;
		12'd 1250 : data_o = 23'b 00101100100011110111111 ;
		12'd 1251 : data_o = 23'b 00101100011100101011011 ;
		12'd 1252 : data_o = 23'b 00101100010101011111010 ;
		12'd 1253 : data_o = 23'b 00101100001110010011011 ;
		12'd 1254 : data_o = 23'b 00101100000111000111101 ;
		12'd 1255 : data_o = 23'b 00101011111111111100010 ;
		12'd 1256 : data_o = 23'b 00101011111000110001001 ;
		12'd 1257 : data_o = 23'b 00101011110001100110010 ;
		12'd 1258 : data_o = 23'b 00101011101010011011101 ;
		12'd 1259 : data_o = 23'b 00101011100011010001010 ;
		12'd 1260 : data_o = 23'b 00101011011100000111001 ;
		12'd 1261 : data_o = 23'b 00101011010100111101010 ;
		12'd 1262 : data_o = 23'b 00101011001101110011101 ;
		12'd 1263 : data_o = 23'b 00101011000110101010010 ;
		12'd 1264 : data_o = 23'b 00101010111111100001001 ;
		12'd 1265 : data_o = 23'b 00101010111000011000011 ;
		12'd 1266 : data_o = 23'b 00101010110001001111110 ;
		12'd 1267 : data_o = 23'b 00101010101010000111011 ;
		12'd 1268 : data_o = 23'b 00101010100010111111011 ;
		12'd 1269 : data_o = 23'b 00101010011011110111100 ;
		12'd 1270 : data_o = 23'b 00101010010100110000000 ;
		12'd 1271 : data_o = 23'b 00101010001101101000101 ;
		12'd 1272 : data_o = 23'b 00101010000110100001101 ;
		12'd 1273 : data_o = 23'b 00101001111111011010110 ;
		12'd 1274 : data_o = 23'b 00101001111000010100010 ;
		12'd 1275 : data_o = 23'b 00101001110001001110000 ;
		12'd 1276 : data_o = 23'b 00101001101010000111111 ;
		12'd 1277 : data_o = 23'b 00101001100011000010001 ;
		12'd 1278 : data_o = 23'b 00101001011011111100101 ;
		12'd 1279 : data_o = 23'b 00101001010100110111011 ;
		12'd 1280 : data_o = 23'b 00101001001101110010010 ;
		12'd 1281 : data_o = 23'b 00101001000110101101100 ;
		12'd 1282 : data_o = 23'b 00101000111111101001000 ;
		12'd 1283 : data_o = 23'b 00101000111000100100110 ;
		12'd 1284 : data_o = 23'b 00101000110001100000110 ;
		12'd 1285 : data_o = 23'b 00101000101010011101000 ;
		12'd 1286 : data_o = 23'b 00101000100011011001100 ;
		12'd 1287 : data_o = 23'b 00101000011100010110001 ;
		12'd 1288 : data_o = 23'b 00101000010101010011001 ;
		12'd 1289 : data_o = 23'b 00101000001110010000011 ;
		12'd 1290 : data_o = 23'b 00101000000111001101111 ;
		12'd 1291 : data_o = 23'b 00101000000000001011101 ;
		12'd 1292 : data_o = 23'b 00100111111001001001101 ;
		12'd 1293 : data_o = 23'b 00100111110010000111111 ;
		12'd 1294 : data_o = 23'b 00100111101011000110011 ;
		12'd 1295 : data_o = 23'b 00100111100100000101001 ;
		12'd 1296 : data_o = 23'b 00100111011101000100001 ;
		12'd 1297 : data_o = 23'b 00100111010110000011011 ;
		12'd 1298 : data_o = 23'b 00100111001111000010111 ;
		12'd 1299 : data_o = 23'b 00100111001000000010101 ;
		12'd 1300 : data_o = 23'b 00100111000001000010101 ;
		12'd 1301 : data_o = 23'b 00100110111010000010111 ;
		12'd 1302 : data_o = 23'b 00100110110011000011011 ;
		12'd 1303 : data_o = 23'b 00100110101100000100001 ;
		12'd 1304 : data_o = 23'b 00100110100101000101000 ;
		12'd 1305 : data_o = 23'b 00100110011110000110010 ;
		12'd 1306 : data_o = 23'b 00100110010111000111110 ;
		12'd 1307 : data_o = 23'b 00100110010000001001100 ;
		12'd 1308 : data_o = 23'b 00100110001001001011100 ;
		12'd 1309 : data_o = 23'b 00100110000010001101110 ;
		12'd 1310 : data_o = 23'b 00100101111011010000010 ;
		12'd 1311 : data_o = 23'b 00100101110100010010111 ;
		12'd 1312 : data_o = 23'b 00100101101101010101111 ;
		12'd 1313 : data_o = 23'b 00100101100110011001001 ;
		12'd 1314 : data_o = 23'b 00100101011111011100101 ;
		12'd 1315 : data_o = 23'b 00100101011000100000010 ;
		12'd 1316 : data_o = 23'b 00100101010001100100010 ;
		12'd 1317 : data_o = 23'b 00100101001010101000011 ;
		12'd 1318 : data_o = 23'b 00100101000011101100111 ;
		12'd 1319 : data_o = 23'b 00100100111100110001101 ;
		12'd 1320 : data_o = 23'b 00100100110101110110100 ;
		12'd 1321 : data_o = 23'b 00100100101110111011110 ;
		12'd 1322 : data_o = 23'b 00100100101000000001001 ;
		12'd 1323 : data_o = 23'b 00100100100001000110110 ;
		12'd 1324 : data_o = 23'b 00100100011010001100110 ;
		12'd 1325 : data_o = 23'b 00100100010011010010111 ;
		12'd 1326 : data_o = 23'b 00100100001100011001010 ;
		12'd 1327 : data_o = 23'b 00100100000101011111111 ;
		12'd 1328 : data_o = 23'b 00100011111110100110111 ;
		12'd 1329 : data_o = 23'b 00100011110111101110000 ;
		12'd 1330 : data_o = 23'b 00100011110000110101011 ;
		12'd 1331 : data_o = 23'b 00100011101001111101000 ;
		12'd 1332 : data_o = 23'b 00100011100011000100111 ;
		12'd 1333 : data_o = 23'b 00100011011100001101000 ;
		12'd 1334 : data_o = 23'b 00100011010101010101011 ;
		12'd 1335 : data_o = 23'b 00100011001110011101111 ;
		12'd 1336 : data_o = 23'b 00100011000111100110110 ;
		12'd 1337 : data_o = 23'b 00100011000000101111111 ;
		12'd 1338 : data_o = 23'b 00100010111001111001001 ;
		12'd 1339 : data_o = 23'b 00100010110011000010110 ;
		12'd 1340 : data_o = 23'b 00100010101100001100100 ;
		12'd 1341 : data_o = 23'b 00100010100101010110101 ;
		12'd 1342 : data_o = 23'b 00100010011110100000111 ;
		12'd 1343 : data_o = 23'b 00100010010111101011100 ;
		12'd 1344 : data_o = 23'b 00100010010000110110010 ;
		12'd 1345 : data_o = 23'b 00100010001010000001010 ;
		12'd 1346 : data_o = 23'b 00100010000011001100100 ;
		12'd 1347 : data_o = 23'b 00100001111100011000000 ;
		12'd 1348 : data_o = 23'b 00100001110101100011110 ;
		12'd 1349 : data_o = 23'b 00100001101110101111110 ;
		12'd 1350 : data_o = 23'b 00100001100111111100000 ;
		12'd 1351 : data_o = 23'b 00100001100001001000011 ;
		12'd 1352 : data_o = 23'b 00100001011010010101001 ;
		12'd 1353 : data_o = 23'b 00100001010011100010000 ;
		12'd 1354 : data_o = 23'b 00100001001100101111010 ;
		12'd 1355 : data_o = 23'b 00100001000101111100101 ;
		12'd 1356 : data_o = 23'b 00100000111111001010010 ;
		12'd 1357 : data_o = 23'b 00100000111000011000010 ;
		12'd 1358 : data_o = 23'b 00100000110001100110011 ;
		12'd 1359 : data_o = 23'b 00100000101010110100110 ;
		12'd 1360 : data_o = 23'b 00100000100100000011011 ;
		12'd 1361 : data_o = 23'b 00100000011101010010001 ;
		12'd 1362 : data_o = 23'b 00100000010110100001010 ;
		12'd 1363 : data_o = 23'b 00100000001111110000101 ;
		12'd 1364 : data_o = 23'b 00100000001001000000001 ;
		12'd 1365 : data_o = 23'b 00100000000010010000000 ;
		12'd 1366 : data_o = 23'b 00011111111011100000000 ;
		12'd 1367 : data_o = 23'b 00011111110100110000010 ;
		12'd 1368 : data_o = 23'b 00011111101110000000110 ;
		12'd 1369 : data_o = 23'b 00011111100111010001100 ;
		12'd 1370 : data_o = 23'b 00011111100000100010100 ;
		12'd 1371 : data_o = 23'b 00011111011001110011110 ;
		12'd 1372 : data_o = 23'b 00011111010011000101010 ;
		12'd 1373 : data_o = 23'b 00011111001100010110111 ;
		12'd 1374 : data_o = 23'b 00011111000101101000111 ;
		12'd 1375 : data_o = 23'b 00011110111110111011000 ;
		12'd 1376 : data_o = 23'b 00011110111000001101011 ;
		12'd 1377 : data_o = 23'b 00011110110001100000000 ;
		12'd 1378 : data_o = 23'b 00011110101010110010111 ;
		12'd 1379 : data_o = 23'b 00011110100100000110000 ;
		12'd 1380 : data_o = 23'b 00011110011101011001011 ;
		12'd 1381 : data_o = 23'b 00011110010110101101000 ;
		12'd 1382 : data_o = 23'b 00011110010000000000110 ;
		12'd 1383 : data_o = 23'b 00011110001001010100110 ;
		12'd 1384 : data_o = 23'b 00011110000010101001001 ;
		12'd 1385 : data_o = 23'b 00011101111011111101101 ;
		12'd 1386 : data_o = 23'b 00011101110101010010011 ;
		12'd 1387 : data_o = 23'b 00011101101110100111011 ;
		12'd 1388 : data_o = 23'b 00011101100111111100101 ;
		12'd 1389 : data_o = 23'b 00011101100001010010000 ;
		12'd 1390 : data_o = 23'b 00011101011010100111110 ;
		12'd 1391 : data_o = 23'b 00011101010011111101101 ;
		12'd 1392 : data_o = 23'b 00011101001101010011110 ;
		12'd 1393 : data_o = 23'b 00011101000110101010001 ;
		12'd 1394 : data_o = 23'b 00011101000000000000110 ;
		12'd 1395 : data_o = 23'b 00011100111001010111101 ;
		12'd 1396 : data_o = 23'b 00011100110010101110110 ;
		12'd 1397 : data_o = 23'b 00011100101100000110000 ;
		12'd 1398 : data_o = 23'b 00011100100101011101100 ;
		12'd 1399 : data_o = 23'b 00011100011110110101011 ;
		12'd 1400 : data_o = 23'b 00011100011000001101011 ;
		12'd 1401 : data_o = 23'b 00011100010001100101101 ;
		12'd 1402 : data_o = 23'b 00011100001010111110000 ;
		12'd 1403 : data_o = 23'b 00011100000100010110110 ;
		12'd 1404 : data_o = 23'b 00011011111101101111101 ;
		12'd 1405 : data_o = 23'b 00011011110111001000111 ;
		12'd 1406 : data_o = 23'b 00011011110000100010010 ;
		12'd 1407 : data_o = 23'b 00011011101001111011111 ;
		12'd 1408 : data_o = 23'b 00011011100011010101110 ;
		12'd 1409 : data_o = 23'b 00011011011100101111110 ;
		12'd 1410 : data_o = 23'b 00011011010110001010001 ;
		12'd 1411 : data_o = 23'b 00011011001111100100101 ;
		12'd 1412 : data_o = 23'b 00011011001000111111011 ;
		12'd 1413 : data_o = 23'b 00011011000010011010011 ;
		12'd 1414 : data_o = 23'b 00011010111011110101101 ;
		12'd 1415 : data_o = 23'b 00011010110101010001001 ;
		12'd 1416 : data_o = 23'b 00011010101110101100110 ;
		12'd 1417 : data_o = 23'b 00011010101000001000110 ;
		12'd 1418 : data_o = 23'b 00011010100001100100111 ;
		12'd 1419 : data_o = 23'b 00011010011011000001010 ;
		12'd 1420 : data_o = 23'b 00011010010100011101111 ;
		12'd 1421 : data_o = 23'b 00011010001101111010101 ;
		12'd 1422 : data_o = 23'b 00011010000111010111110 ;
		12'd 1423 : data_o = 23'b 00011010000000110101000 ;
		12'd 1424 : data_o = 23'b 00011001111010010010100 ;
		12'd 1425 : data_o = 23'b 00011001110011110000010 ;
		12'd 1426 : data_o = 23'b 00011001101101001110010 ;
		12'd 1427 : data_o = 23'b 00011001100110101100100 ;
		12'd 1428 : data_o = 23'b 00011001100000001010111 ;
		12'd 1429 : data_o = 23'b 00011001011001101001100 ;
		12'd 1430 : data_o = 23'b 00011001010011001000011 ;
		12'd 1431 : data_o = 23'b 00011001001100100111100 ;
		12'd 1432 : data_o = 23'b 00011001000110000110111 ;
		12'd 1433 : data_o = 23'b 00011000111111100110011 ;
		12'd 1434 : data_o = 23'b 00011000111001000110001 ;
		12'd 1435 : data_o = 23'b 00011000110010100110001 ;
		12'd 1436 : data_o = 23'b 00011000101100000110011 ;
		12'd 1437 : data_o = 23'b 00011000100101100110111 ;
		12'd 1438 : data_o = 23'b 00011000011111000111100 ;
		12'd 1439 : data_o = 23'b 00011000011000101000100 ;
		12'd 1440 : data_o = 23'b 00011000010010001001101 ;
		12'd 1441 : data_o = 23'b 00011000001011101011000 ;
		12'd 1442 : data_o = 23'b 00011000000101001100100 ;
		12'd 1443 : data_o = 23'b 00010111111110101110011 ;
		12'd 1444 : data_o = 23'b 00010111111000010000011 ;
		12'd 1445 : data_o = 23'b 00010111110001110010101 ;
		12'd 1446 : data_o = 23'b 00010111101011010101001 ;
		12'd 1447 : data_o = 23'b 00010111100100110111110 ;
		12'd 1448 : data_o = 23'b 00010111011110011010110 ;
		12'd 1449 : data_o = 23'b 00010111010111111101111 ;
		12'd 1450 : data_o = 23'b 00010111010001100001010 ;
		12'd 1451 : data_o = 23'b 00010111001011000100111 ;
		12'd 1452 : data_o = 23'b 00010111000100101000101 ;
		12'd 1453 : data_o = 23'b 00010110111110001100110 ;
		12'd 1454 : data_o = 23'b 00010110110111110001000 ;
		12'd 1455 : data_o = 23'b 00010110110001010101100 ;
		12'd 1456 : data_o = 23'b 00010110101010111010001 ;
		12'd 1457 : data_o = 23'b 00010110100100011111001 ;
		12'd 1458 : data_o = 23'b 00010110011110000100010 ;
		12'd 1459 : data_o = 23'b 00010110010111101001101 ;
		12'd 1460 : data_o = 23'b 00010110010001001111010 ;
		12'd 1461 : data_o = 23'b 00010110001010110101000 ;
		12'd 1462 : data_o = 23'b 00010110000100011011001 ;
		12'd 1463 : data_o = 23'b 00010101111110000001011 ;
		12'd 1464 : data_o = 23'b 00010101110111100111111 ;
		12'd 1465 : data_o = 23'b 00010101110001001110100 ;
		12'd 1466 : data_o = 23'b 00010101101010110101100 ;
		12'd 1467 : data_o = 23'b 00010101100100011100101 ;
		12'd 1468 : data_o = 23'b 00010101011110000100000 ;
		12'd 1469 : data_o = 23'b 00010101010111101011100 ;
		12'd 1470 : data_o = 23'b 00010101010001010011011 ;
		12'd 1471 : data_o = 23'b 00010101001010111011011 ;
		12'd 1472 : data_o = 23'b 00010101000100100011101 ;
		12'd 1473 : data_o = 23'b 00010100111110001100001 ;
		12'd 1474 : data_o = 23'b 00010100110111110100110 ;
		12'd 1475 : data_o = 23'b 00010100110001011101101 ;
		12'd 1476 : data_o = 23'b 00010100101011000110110 ;
		12'd 1477 : data_o = 23'b 00010100100100110000001 ;
		12'd 1478 : data_o = 23'b 00010100011110011001110 ;
		12'd 1479 : data_o = 23'b 00010100011000000011100 ;
		12'd 1480 : data_o = 23'b 00010100010001101101100 ;
		12'd 1481 : data_o = 23'b 00010100001011010111110 ;
		12'd 1482 : data_o = 23'b 00010100000101000010001 ;
		12'd 1483 : data_o = 23'b 00010011111110101100110 ;
		12'd 1484 : data_o = 23'b 00010011111000010111101 ;
		12'd 1485 : data_o = 23'b 00010011110010000010110 ;
		12'd 1486 : data_o = 23'b 00010011101011101110000 ;
		12'd 1487 : data_o = 23'b 00010011100101011001101 ;
		12'd 1488 : data_o = 23'b 00010011011111000101010 ;
		12'd 1489 : data_o = 23'b 00010011011000110001010 ;
		12'd 1490 : data_o = 23'b 00010011010010011101100 ;
		12'd 1491 : data_o = 23'b 00010011001100001001111 ;
		12'd 1492 : data_o = 23'b 00010011000101110110100 ;
		12'd 1493 : data_o = 23'b 00010010111111100011010 ;
		12'd 1494 : data_o = 23'b 00010010111001010000010 ;
		12'd 1495 : data_o = 23'b 00010010110010111101100 ;
		12'd 1496 : data_o = 23'b 00010010101100101011000 ;
		12'd 1497 : data_o = 23'b 00010010100110011000110 ;
		12'd 1498 : data_o = 23'b 00010010100000000110101 ;
		12'd 1499 : data_o = 23'b 00010010011001110100110 ;
		12'd 1500 : data_o = 23'b 00010010010011100011001 ;
		12'd 1501 : data_o = 23'b 00010010001101010001101 ;
		12'd 1502 : data_o = 23'b 00010010000111000000011 ;
		12'd 1503 : data_o = 23'b 00010010000000101111011 ;
		12'd 1504 : data_o = 23'b 00010001111010011110101 ;
		12'd 1505 : data_o = 23'b 00010001110100001110000 ;
		12'd 1506 : data_o = 23'b 00010001101101111101101 ;
		12'd 1507 : data_o = 23'b 00010001100111101101100 ;
		12'd 1508 : data_o = 23'b 00010001100001011101100 ;
		12'd 1509 : data_o = 23'b 00010001011011001101110 ;
		12'd 1510 : data_o = 23'b 00010001010100111110010 ;
		12'd 1511 : data_o = 23'b 00010001001110101111000 ;
		12'd 1512 : data_o = 23'b 00010001001000011111111 ;
		12'd 1513 : data_o = 23'b 00010001000010010001000 ;
		12'd 1514 : data_o = 23'b 00010000111100000010011 ;
		12'd 1515 : data_o = 23'b 00010000110101110011111 ;
		12'd 1516 : data_o = 23'b 00010000101111100101101 ;
		12'd 1517 : data_o = 23'b 00010000101001010111101 ;
		12'd 1518 : data_o = 23'b 00010000100011001001110 ;
		12'd 1519 : data_o = 23'b 00010000011100111100010 ;
		12'd 1520 : data_o = 23'b 00010000010110101110110 ;
		12'd 1521 : data_o = 23'b 00010000010000100001101 ;
		12'd 1522 : data_o = 23'b 00010000001010010100101 ;
		12'd 1523 : data_o = 23'b 00010000000100000111111 ;
		12'd 1524 : data_o = 23'b 00001111111101111011011 ;
		12'd 1525 : data_o = 23'b 00001111110111101111000 ;
		12'd 1526 : data_o = 23'b 00001111110001100010111 ;
		12'd 1527 : data_o = 23'b 00001111101011010111000 ;
		12'd 1528 : data_o = 23'b 00001111100101001011011 ;
		12'd 1529 : data_o = 23'b 00001111011110111111111 ;
		12'd 1530 : data_o = 23'b 00001111011000110100101 ;
		12'd 1531 : data_o = 23'b 00001111010010101001100 ;
		12'd 1532 : data_o = 23'b 00001111001100011110101 ;
		12'd 1533 : data_o = 23'b 00001111000110010100000 ;
		12'd 1534 : data_o = 23'b 00001111000000001001101 ;
		12'd 1535 : data_o = 23'b 00001110111001111111011 ;
		12'd 1536 : data_o = 23'b 00001110110011110101011 ;
		12'd 1537 : data_o = 23'b 00001110101101101011100 ;
		12'd 1538 : data_o = 23'b 00001110100111100010000 ;
		12'd 1539 : data_o = 23'b 00001110100001011000101 ;
		12'd 1540 : data_o = 23'b 00001110011011001111011 ;
		12'd 1541 : data_o = 23'b 00001110010101000110100 ;
		12'd 1542 : data_o = 23'b 00001110001110111101110 ;
		12'd 1543 : data_o = 23'b 00001110001000110101001 ;
		12'd 1544 : data_o = 23'b 00001110000010101100111 ;
		12'd 1545 : data_o = 23'b 00001101111100100100110 ;
		12'd 1546 : data_o = 23'b 00001101110110011100110 ;
		12'd 1547 : data_o = 23'b 00001101110000010101000 ;
		12'd 1548 : data_o = 23'b 00001101101010001101100 ;
		12'd 1549 : data_o = 23'b 00001101100100000110010 ;
		12'd 1550 : data_o = 23'b 00001101011101111111001 ;
		12'd 1551 : data_o = 23'b 00001101010111111000010 ;
		12'd 1552 : data_o = 23'b 00001101010001110001101 ;
		12'd 1553 : data_o = 23'b 00001101001011101011001 ;
		12'd 1554 : data_o = 23'b 00001101000101100100111 ;
		12'd 1555 : data_o = 23'b 00001100111111011110111 ;
		12'd 1556 : data_o = 23'b 00001100111001011001000 ;
		12'd 1557 : data_o = 23'b 00001100110011010011011 ;
		12'd 1558 : data_o = 23'b 00001100101101001110000 ;
		12'd 1559 : data_o = 23'b 00001100100111001000110 ;
		12'd 1560 : data_o = 23'b 00001100100001000011110 ;
		12'd 1561 : data_o = 23'b 00001100011010111110111 ;
		12'd 1562 : data_o = 23'b 00001100010100111010010 ;
		12'd 1563 : data_o = 23'b 00001100001110110101111 ;
		12'd 1564 : data_o = 23'b 00001100001000110001110 ;
		12'd 1565 : data_o = 23'b 00001100000010101101110 ;
		12'd 1566 : data_o = 23'b 00001011111100101010000 ;
		12'd 1567 : data_o = 23'b 00001011110110100110011 ;
		12'd 1568 : data_o = 23'b 00001011110000100011000 ;
		12'd 1569 : data_o = 23'b 00001011101010011111111 ;
		12'd 1570 : data_o = 23'b 00001011100100011100111 ;
		12'd 1571 : data_o = 23'b 00001011011110011010001 ;
		12'd 1572 : data_o = 23'b 00001011011000010111101 ;
		12'd 1573 : data_o = 23'b 00001011010010010101010 ;
		12'd 1574 : data_o = 23'b 00001011001100010011001 ;
		12'd 1575 : data_o = 23'b 00001011000110010001001 ;
		12'd 1576 : data_o = 23'b 00001011000000001111011 ;
		12'd 1577 : data_o = 23'b 00001010111010001101111 ;
		12'd 1578 : data_o = 23'b 00001010110100001100101 ;
		12'd 1579 : data_o = 23'b 00001010101110001011100 ;
		12'd 1580 : data_o = 23'b 00001010101000001010100 ;
		12'd 1581 : data_o = 23'b 00001010100010001001111 ;
		12'd 1582 : data_o = 23'b 00001010011100001001010 ;
		12'd 1583 : data_o = 23'b 00001010010110001001000 ;
		12'd 1584 : data_o = 23'b 00001010010000001000111 ;
		12'd 1585 : data_o = 23'b 00001010001010001001000 ;
		12'd 1586 : data_o = 23'b 00001010000100001001010 ;
		12'd 1587 : data_o = 23'b 00001001111110001001110 ;
		12'd 1588 : data_o = 23'b 00001001111000001010100 ;
		12'd 1589 : data_o = 23'b 00001001110010001011011 ;
		12'd 1590 : data_o = 23'b 00001001101100001100100 ;
		12'd 1591 : data_o = 23'b 00001001100110001101111 ;
		12'd 1592 : data_o = 23'b 00001001100000001111011 ;
		12'd 1593 : data_o = 23'b 00001001011010010001001 ;
		12'd 1594 : data_o = 23'b 00001001010100010011000 ;
		12'd 1595 : data_o = 23'b 00001001001110010101001 ;
		12'd 1596 : data_o = 23'b 00001001001000010111011 ;
		12'd 1597 : data_o = 23'b 00001001000010011010000 ;
		12'd 1598 : data_o = 23'b 00001000111100011100101 ;
		12'd 1599 : data_o = 23'b 00001000110110011111101 ;
		12'd 1600 : data_o = 23'b 00001000110000100010110 ;
		12'd 1601 : data_o = 23'b 00001000101010100110000 ;
		12'd 1602 : data_o = 23'b 00001000100100101001100 ;
		12'd 1603 : data_o = 23'b 00001000011110101101010 ;
		12'd 1604 : data_o = 23'b 00001000011000110001010 ;
		12'd 1605 : data_o = 23'b 00001000010010110101011 ;
		12'd 1606 : data_o = 23'b 00001000001100111001101 ;
		12'd 1607 : data_o = 23'b 00001000000110111110001 ;
		12'd 1608 : data_o = 23'b 00001000000001000010111 ;
		12'd 1609 : data_o = 23'b 00000111111011000111111 ;
		12'd 1610 : data_o = 23'b 00000111110101001101000 ;
		12'd 1611 : data_o = 23'b 00000111101111010010010 ;
		12'd 1612 : data_o = 23'b 00000111101001010111110 ;
		12'd 1613 : data_o = 23'b 00000111100011011101100 ;
		12'd 1614 : data_o = 23'b 00000111011101100011011 ;
		12'd 1615 : data_o = 23'b 00000111010111101001100 ;
		12'd 1616 : data_o = 23'b 00000111010001101111111 ;
		12'd 1617 : data_o = 23'b 00000111001011110110011 ;
		12'd 1618 : data_o = 23'b 00000111000101111101001 ;
		12'd 1619 : data_o = 23'b 00000111000000000100000 ;
		12'd 1620 : data_o = 23'b 00000110111010001011001 ;
		12'd 1621 : data_o = 23'b 00000110110100010010011 ;
		12'd 1622 : data_o = 23'b 00000110101110011001111 ;
		12'd 1623 : data_o = 23'b 00000110101000100001101 ;
		12'd 1624 : data_o = 23'b 00000110100010101001100 ;
		12'd 1625 : data_o = 23'b 00000110011100110001101 ;
		12'd 1626 : data_o = 23'b 00000110010110111001111 ;
		12'd 1627 : data_o = 23'b 00000110010001000010011 ;
		12'd 1628 : data_o = 23'b 00000110001011001011001 ;
		12'd 1629 : data_o = 23'b 00000110000101010100000 ;
		12'd 1630 : data_o = 23'b 00000101111111011101000 ;
		12'd 1631 : data_o = 23'b 00000101111001100110011 ;
		12'd 1632 : data_o = 23'b 00000101110011101111110 ;
		12'd 1633 : data_o = 23'b 00000101101101111001100 ;
		12'd 1634 : data_o = 23'b 00000101101000000011011 ;
		12'd 1635 : data_o = 23'b 00000101100010001101011 ;
		12'd 1636 : data_o = 23'b 00000101011100010111101 ;
		12'd 1637 : data_o = 23'b 00000101010110100010001 ;
		12'd 1638 : data_o = 23'b 00000101010000101100110 ;
		12'd 1639 : data_o = 23'b 00000101001010110111101 ;
		12'd 1640 : data_o = 23'b 00000101000101000010101 ;
		12'd 1641 : data_o = 23'b 00000100111111001101111 ;
		12'd 1642 : data_o = 23'b 00000100111001011001010 ;
		12'd 1643 : data_o = 23'b 00000100110011100100111 ;
		12'd 1644 : data_o = 23'b 00000100101101110000110 ;
		12'd 1645 : data_o = 23'b 00000100100111111100110 ;
		12'd 1646 : data_o = 23'b 00000100100010001000111 ;
		12'd 1647 : data_o = 23'b 00000100011100010101011 ;
		12'd 1648 : data_o = 23'b 00000100010110100001111 ;
		12'd 1649 : data_o = 23'b 00000100010000101110110 ;
		12'd 1650 : data_o = 23'b 00000100001010111011101 ;
		12'd 1651 : data_o = 23'b 00000100000101001000111 ;
		12'd 1652 : data_o = 23'b 00000011111111010110010 ;
		12'd 1653 : data_o = 23'b 00000011111001100011110 ;
		12'd 1654 : data_o = 23'b 00000011110011110001100 ;
		12'd 1655 : data_o = 23'b 00000011101101111111100 ;
		12'd 1656 : data_o = 23'b 00000011101000001101101 ;
		12'd 1657 : data_o = 23'b 00000011100010011100000 ;
		12'd 1658 : data_o = 23'b 00000011011100101010100 ;
		12'd 1659 : data_o = 23'b 00000011010110111001010 ;
		12'd 1660 : data_o = 23'b 00000011010001001000001 ;
		12'd 1661 : data_o = 23'b 00000011001011010111010 ;
		12'd 1662 : data_o = 23'b 00000011000101100110100 ;
		12'd 1663 : data_o = 23'b 00000010111111110110000 ;
		12'd 1664 : data_o = 23'b 00000010111010000101110 ;
		12'd 1665 : data_o = 23'b 00000010110100010101100 ;
		12'd 1666 : data_o = 23'b 00000010101110100101101 ;
		12'd 1667 : data_o = 23'b 00000010101000110101111 ;
		12'd 1668 : data_o = 23'b 00000010100011000110011 ;
		12'd 1669 : data_o = 23'b 00000010011101010111000 ;
		12'd 1670 : data_o = 23'b 00000010010111100111110 ;
		12'd 1671 : data_o = 23'b 00000010010001111000110 ;
		12'd 1672 : data_o = 23'b 00000010001100001010000 ;
		12'd 1673 : data_o = 23'b 00000010000110011011011 ;
		12'd 1674 : data_o = 23'b 00000010000000101101000 ;
		12'd 1675 : data_o = 23'b 00000001111010111110110 ;
		12'd 1676 : data_o = 23'b 00000001110101010000110 ;
		12'd 1677 : data_o = 23'b 00000001101111100010111 ;
		12'd 1678 : data_o = 23'b 00000001101001110101010 ;
		12'd 1679 : data_o = 23'b 00000001100100000111111 ;
		12'd 1680 : data_o = 23'b 00000001011110011010100 ;
		12'd 1681 : data_o = 23'b 00000001011000101101100 ;
		12'd 1682 : data_o = 23'b 00000001010011000000101 ;
		12'd 1683 : data_o = 23'b 00000001001101010011111 ;
		12'd 1684 : data_o = 23'b 00000001000111100111011 ;
		12'd 1685 : data_o = 23'b 00000001000001111011001 ;
		12'd 1686 : data_o = 23'b 00000000111100001110111 ;
		12'd 1687 : data_o = 23'b 00000000110110100011000 ;
		12'd 1688 : data_o = 23'b 00000000110000110111010 ;
		12'd 1689 : data_o = 23'b 00000000101011001011101 ;
		12'd 1690 : data_o = 23'b 00000000100101100000010 ;
		12'd 1691 : data_o = 23'b 00000000011111110101001 ;
		12'd 1692 : data_o = 23'b 00000000011010001010001 ;
		12'd 1693 : data_o = 23'b 00000000010100011111010 ;
		12'd 1694 : data_o = 23'b 00000000001110110100101 ;
		12'd 1695 : data_o = 23'b 00000000001001001010010 ;
		12'd 1696 : data_o = 23'b 00000000000011100000000 ;
		12'd 1697 : data_o = 23'b 11111111111011101011111 ;
		12'd 1698 : data_o = 23'b 11111111110000011000001 ;
		12'd 1699 : data_o = 23'b 11111111100101000100110 ;
		12'd 1700 : data_o = 23'b 11111111011001110001110 ;
		12'd 1701 : data_o = 23'b 11111111001110011111001 ;
		12'd 1702 : data_o = 23'b 11111111000011001100111 ;
		12'd 1703 : data_o = 23'b 11111110110111111011000 ;
		12'd 1704 : data_o = 23'b 11111110101100101001100 ;
		12'd 1705 : data_o = 23'b 11111110100001011000011 ;
		12'd 1706 : data_o = 23'b 11111110010110000111101 ;
		12'd 1707 : data_o = 23'b 11111110001010110111010 ;
		12'd 1708 : data_o = 23'b 11111101111111100111010 ;
		12'd 1709 : data_o = 23'b 11111101110100010111101 ;
		12'd 1710 : data_o = 23'b 11111101101001001000011 ;
		12'd 1711 : data_o = 23'b 11111101011101111001100 ;
		12'd 1712 : data_o = 23'b 11111101010010101010111 ;
		12'd 1713 : data_o = 23'b 11111101000111011100110 ;
		12'd 1714 : data_o = 23'b 11111100111100001111000 ;
		12'd 1715 : data_o = 23'b 11111100110001000001101 ;
		12'd 1716 : data_o = 23'b 11111100100101110100100 ;
		12'd 1717 : data_o = 23'b 11111100011010100111111 ;
		12'd 1718 : data_o = 23'b 11111100001111011011100 ;
		12'd 1719 : data_o = 23'b 11111100000100001111101 ;
		12'd 1720 : data_o = 23'b 11111011111001000100000 ;
		12'd 1721 : data_o = 23'b 11111011101101111000111 ;
		12'd 1722 : data_o = 23'b 11111011100010101110000 ;
		12'd 1723 : data_o = 23'b 11111011010111100011101 ;
		12'd 1724 : data_o = 23'b 11111011001100011001100 ;
		12'd 1725 : data_o = 23'b 11111011000001001111110 ;
		12'd 1726 : data_o = 23'b 11111010110110000110011 ;
		12'd 1727 : data_o = 23'b 11111010101010111101011 ;
		12'd 1728 : data_o = 23'b 11111010011111110100110 ;
		12'd 1729 : data_o = 23'b 11111010010100101100100 ;
		12'd 1730 : data_o = 23'b 11111010001001100100101 ;
		12'd 1731 : data_o = 23'b 11111001111110011101001 ;
		12'd 1732 : data_o = 23'b 11111001110011010110000 ;
		12'd 1733 : data_o = 23'b 11111001101000001111010 ;
		12'd 1734 : data_o = 23'b 11111001011101001000110 ;
		12'd 1735 : data_o = 23'b 11111001010010000010110 ;
		12'd 1736 : data_o = 23'b 11111001000110111101000 ;
		12'd 1737 : data_o = 23'b 11111000111011110111110 ;
		12'd 1738 : data_o = 23'b 11111000110000110010110 ;
		12'd 1739 : data_o = 23'b 11111000100101101110001 ;
		12'd 1740 : data_o = 23'b 11111000011010101001111 ;
		12'd 1741 : data_o = 23'b 11111000001111100110000 ;
		12'd 1742 : data_o = 23'b 11111000000100100010100 ;
		12'd 1743 : data_o = 23'b 11110111111001011111011 ;
		12'd 1744 : data_o = 23'b 11110111101110011100101 ;
		12'd 1745 : data_o = 23'b 11110111100011011010010 ;
		12'd 1746 : data_o = 23'b 11110111011000011000001 ;
		12'd 1747 : data_o = 23'b 11110111001101010110100 ;
		12'd 1748 : data_o = 23'b 11110111000010010101001 ;
		12'd 1749 : data_o = 23'b 11110110110111010100010 ;
		12'd 1750 : data_o = 23'b 11110110101100010011101 ;
		12'd 1751 : data_o = 23'b 11110110100001010011011 ;
		12'd 1752 : data_o = 23'b 11110110010110010011100 ;
		12'd 1753 : data_o = 23'b 11110110001011010100000 ;
		12'd 1754 : data_o = 23'b 11110110000000010100110 ;
		12'd 1755 : data_o = 23'b 11110101110101010110000 ;
		12'd 1756 : data_o = 23'b 11110101101010010111100 ;
		12'd 1757 : data_o = 23'b 11110101011111011001100 ;
		12'd 1758 : data_o = 23'b 11110101010100011011110 ;
		12'd 1759 : data_o = 23'b 11110101001001011110011 ;
		12'd 1760 : data_o = 23'b 11110100111110100001011 ;
		12'd 1761 : data_o = 23'b 11110100110011100100110 ;
		12'd 1762 : data_o = 23'b 11110100101000101000100 ;
		12'd 1763 : data_o = 23'b 11110100011101101100100 ;
		12'd 1764 : data_o = 23'b 11110100010010110001000 ;
		12'd 1765 : data_o = 23'b 11110100000111110101110 ;
		12'd 1766 : data_o = 23'b 11110011111100111010111 ;
		12'd 1767 : data_o = 23'b 11110011110010000000011 ;
		12'd 1768 : data_o = 23'b 11110011100111000110010 ;
		12'd 1769 : data_o = 23'b 11110011011100001100100 ;
		12'd 1770 : data_o = 23'b 11110011010001010011001 ;
		12'd 1771 : data_o = 23'b 11110011000110011010000 ;
		12'd 1772 : data_o = 23'b 11110010111011100001011 ;
		12'd 1773 : data_o = 23'b 11110010110000101001000 ;
		12'd 1774 : data_o = 23'b 11110010100101110001000 ;
		12'd 1775 : data_o = 23'b 11110010011010111001011 ;
		12'd 1776 : data_o = 23'b 11110010010000000010000 ;
		12'd 1777 : data_o = 23'b 11110010000101001011001 ;
		12'd 1778 : data_o = 23'b 11110001111010010100100 ;
		12'd 1779 : data_o = 23'b 11110001101111011110011 ;
		12'd 1780 : data_o = 23'b 11110001100100101000100 ;
		12'd 1781 : data_o = 23'b 11110001011001110011000 ;
		12'd 1782 : data_o = 23'b 11110001001110111101110 ;
		12'd 1783 : data_o = 23'b 11110001000100001001000 ;
		12'd 1784 : data_o = 23'b 11110000111001010100100 ;
		12'd 1785 : data_o = 23'b 11110000101110100000100 ;
		12'd 1786 : data_o = 23'b 11110000100011101100110 ;
		12'd 1787 : data_o = 23'b 11110000011000111001011 ;
		12'd 1788 : data_o = 23'b 11110000001110000110010 ;
		12'd 1789 : data_o = 23'b 11110000000011010011101 ;
		12'd 1790 : data_o = 23'b 11101111111000100001010 ;
		12'd 1791 : data_o = 23'b 11101111101101101111010 ;
		12'd 1792 : data_o = 23'b 11101111100010111101101 ;
		12'd 1793 : data_o = 23'b 11101111011000001100011 ;
		12'd 1794 : data_o = 23'b 11101111001101011011011 ;
		12'd 1795 : data_o = 23'b 11101111000010101010111 ;
		12'd 1796 : data_o = 23'b 11101110110111111010101 ;
		12'd 1797 : data_o = 23'b 11101110101101001010110 ;
		12'd 1798 : data_o = 23'b 11101110100010011011010 ;
		12'd 1799 : data_o = 23'b 11101110010111101100000 ;
		12'd 1800 : data_o = 23'b 11101110001100111101010 ;
		12'd 1801 : data_o = 23'b 11101110000010001110110 ;
		12'd 1802 : data_o = 23'b 11101101110111100000101 ;
		12'd 1803 : data_o = 23'b 11101101101100110010111 ;
		12'd 1804 : data_o = 23'b 11101101100010000101011 ;
		12'd 1805 : data_o = 23'b 11101101010111011000010 ;
		12'd 1806 : data_o = 23'b 11101101001100101011101 ;
		12'd 1807 : data_o = 23'b 11101101000001111111010 ;
		12'd 1808 : data_o = 23'b 11101100110111010011001 ;
		12'd 1809 : data_o = 23'b 11101100101100100111100 ;
		12'd 1810 : data_o = 23'b 11101100100001111100001 ;
		12'd 1811 : data_o = 23'b 11101100010111010001001 ;
		12'd 1812 : data_o = 23'b 11101100001100100110100 ;
		12'd 1813 : data_o = 23'b 11101100000001111100001 ;
		12'd 1814 : data_o = 23'b 11101011110111010010010 ;
		12'd 1815 : data_o = 23'b 11101011101100101000101 ;
		12'd 1816 : data_o = 23'b 11101011100001111111011 ;
		12'd 1817 : data_o = 23'b 11101011010111010110011 ;
		12'd 1818 : data_o = 23'b 11101011001100101101111 ;
		12'd 1819 : data_o = 23'b 11101011000010000101101 ;
		12'd 1820 : data_o = 23'b 11101010110111011101110 ;
		12'd 1821 : data_o = 23'b 11101010101100110110001 ;
		12'd 1822 : data_o = 23'b 11101010100010001111000 ;
		12'd 1823 : data_o = 23'b 11101010010111101000001 ;
		12'd 1824 : data_o = 23'b 11101010001101000001101 ;
		12'd 1825 : data_o = 23'b 11101010000010011011100 ;
		12'd 1826 : data_o = 23'b 11101001110111110101101 ;
		12'd 1827 : data_o = 23'b 11101001101101010000001 ;
		12'd 1828 : data_o = 23'b 11101001100010101011000 ;
		12'd 1829 : data_o = 23'b 11101001011000000110010 ;
		12'd 1830 : data_o = 23'b 11101001001101100001110 ;
		12'd 1831 : data_o = 23'b 11101001000010111101101 ;
		12'd 1832 : data_o = 23'b 11101000111000011001111 ;
		12'd 1833 : data_o = 23'b 11101000101101110110100 ;
		12'd 1834 : data_o = 23'b 11101000100011010011011 ;
		12'd 1835 : data_o = 23'b 11101000011000110000101 ;
		12'd 1836 : data_o = 23'b 11101000001110001110010 ;
		12'd 1837 : data_o = 23'b 11101000000011101100010 ;
		12'd 1838 : data_o = 23'b 11100111111001001010100 ;
		12'd 1839 : data_o = 23'b 11100111101110101001001 ;
		12'd 1840 : data_o = 23'b 11100111100100001000001 ;
		12'd 1841 : data_o = 23'b 11100111011001100111011 ;
		12'd 1842 : data_o = 23'b 11100111001111000111000 ;
		12'd 1843 : data_o = 23'b 11100111000100100111000 ;
		12'd 1844 : data_o = 23'b 11100110111010000111011 ;
		12'd 1845 : data_o = 23'b 11100110101111101000000 ;
		12'd 1846 : data_o = 23'b 11100110100101001001000 ;
		12'd 1847 : data_o = 23'b 11100110011010101010011 ;
		12'd 1848 : data_o = 23'b 11100110010000001100000 ;
		12'd 1849 : data_o = 23'b 11100110000101101110000 ;
		12'd 1850 : data_o = 23'b 11100101111011010000011 ;
		12'd 1851 : data_o = 23'b 11100101110000110011001 ;
		12'd 1852 : data_o = 23'b 11100101100110010110001 ;
		12'd 1853 : data_o = 23'b 11100101011011111001100 ;
		12'd 1854 : data_o = 23'b 11100101010001011101010 ;
		12'd 1855 : data_o = 23'b 11100101000111000001010 ;
		12'd 1856 : data_o = 23'b 11100100111100100101101 ;
		12'd 1857 : data_o = 23'b 11100100110010001010011 ;
		12'd 1858 : data_o = 23'b 11100100100111101111011 ;
		12'd 1859 : data_o = 23'b 11100100011101010100110 ;
		12'd 1860 : data_o = 23'b 11100100010010111010100 ;
		12'd 1861 : data_o = 23'b 11100100001000100000100 ;
		12'd 1862 : data_o = 23'b 11100011111110000111000 ;
		12'd 1863 : data_o = 23'b 11100011110011101101101 ;
		12'd 1864 : data_o = 23'b 11100011101001010100110 ;
		12'd 1865 : data_o = 23'b 11100011011110111100001 ;
		12'd 1866 : data_o = 23'b 11100011010100100011111 ;
		12'd 1867 : data_o = 23'b 11100011001010001011111 ;
		12'd 1868 : data_o = 23'b 11100010111111110100011 ;
		12'd 1869 : data_o = 23'b 11100010110101011101001 ;
		12'd 1870 : data_o = 23'b 11100010101011000110001 ;
		12'd 1871 : data_o = 23'b 11100010100000101111100 ;
		12'd 1872 : data_o = 23'b 11100010010110011001010 ;
		12'd 1873 : data_o = 23'b 11100010001100000011011 ;
		12'd 1874 : data_o = 23'b 11100010000001101101110 ;
		12'd 1875 : data_o = 23'b 11100001110111011000100 ;
		12'd 1876 : data_o = 23'b 11100001101101000011100 ;
		12'd 1877 : data_o = 23'b 11100001100010101110111 ;
		12'd 1878 : data_o = 23'b 11100001011000011010101 ;
		12'd 1879 : data_o = 23'b 11100001001110000110110 ;
		12'd 1880 : data_o = 23'b 11100001000011110011001 ;
		12'd 1881 : data_o = 23'b 11100000111001011111111 ;
		12'd 1882 : data_o = 23'b 11100000101111001100111 ;
		12'd 1883 : data_o = 23'b 11100000100100111010010 ;
		12'd 1884 : data_o = 23'b 11100000011010101000000 ;
		12'd 1885 : data_o = 23'b 11100000010000010110000 ;
		12'd 1886 : data_o = 23'b 11100000000110000100011 ;
		12'd 1887 : data_o = 23'b 11011111111011110011001 ;
		12'd 1888 : data_o = 23'b 11011111110001100010001 ;
		12'd 1889 : data_o = 23'b 11011111100111010001100 ;
		12'd 1890 : data_o = 23'b 11011111011101000001001 ;
		12'd 1891 : data_o = 23'b 11011111010010110001010 ;
		12'd 1892 : data_o = 23'b 11011111001000100001100 ;
		12'd 1893 : data_o = 23'b 11011110111110010010010 ;
		12'd 1894 : data_o = 23'b 11011110110100000011010 ;
		12'd 1895 : data_o = 23'b 11011110101001110100100 ;
		12'd 1896 : data_o = 23'b 11011110011111100110010 ;
		12'd 1897 : data_o = 23'b 11011110010101011000010 ;
		12'd 1898 : data_o = 23'b 11011110001011001010100 ;
		12'd 1899 : data_o = 23'b 11011110000000111101001 ;
		12'd 1900 : data_o = 23'b 11011101110110110000001 ;
		12'd 1901 : data_o = 23'b 11011101101100100011011 ;
		12'd 1902 : data_o = 23'b 11011101100010010111000 ;
		12'd 1903 : data_o = 23'b 11011101011000001011000 ;
		12'd 1904 : data_o = 23'b 11011101001101111111010 ;
		12'd 1905 : data_o = 23'b 11011101000011110011111 ;
		12'd 1906 : data_o = 23'b 11011100111001101000110 ;
		12'd 1907 : data_o = 23'b 11011100101111011110000 ;
		12'd 1908 : data_o = 23'b 11011100100101010011101 ;
		12'd 1909 : data_o = 23'b 11011100011011001001100 ;
		12'd 1910 : data_o = 23'b 11011100010000111111110 ;
		12'd 1911 : data_o = 23'b 11011100000110110110010 ;
		12'd 1912 : data_o = 23'b 11011011111100101101001 ;
		12'd 1913 : data_o = 23'b 11011011110010100100011 ;
		12'd 1914 : data_o = 23'b 11011011101000011011111 ;
		12'd 1915 : data_o = 23'b 11011011011110010011110 ;
		12'd 1916 : data_o = 23'b 11011011010100001011111 ;
		12'd 1917 : data_o = 23'b 11011011001010000100011 ;
		12'd 1918 : data_o = 23'b 11011010111111111101010 ;
		12'd 1919 : data_o = 23'b 11011010110101110110011 ;
		12'd 1920 : data_o = 23'b 11011010101011101111111 ;
		12'd 1921 : data_o = 23'b 11011010100001101001101 ;
		12'd 1922 : data_o = 23'b 11011010010111100011110 ;
		12'd 1923 : data_o = 23'b 11011010001101011110001 ;
		12'd 1924 : data_o = 23'b 11011010000011011000111 ;
		12'd 1925 : data_o = 23'b 11011001111001010100000 ;
		12'd 1926 : data_o = 23'b 11011001101111001111011 ;
		12'd 1927 : data_o = 23'b 11011001100101001011001 ;
		12'd 1928 : data_o = 23'b 11011001011011000111001 ;
		12'd 1929 : data_o = 23'b 11011001010001000011100 ;
		12'd 1930 : data_o = 23'b 11011001000111000000001 ;
		12'd 1931 : data_o = 23'b 11011000111100111101001 ;
		12'd 1932 : data_o = 23'b 11011000110010111010100 ;
		12'd 1933 : data_o = 23'b 11011000101000111000001 ;
		12'd 1934 : data_o = 23'b 11011000011110110110000 ;
		12'd 1935 : data_o = 23'b 11011000010100110100010 ;
		12'd 1936 : data_o = 23'b 11011000001010110010111 ;
		12'd 1937 : data_o = 23'b 11011000000000110001110 ;
		12'd 1938 : data_o = 23'b 11010111110110110001000 ;
		12'd 1939 : data_o = 23'b 11010111101100110000101 ;
		12'd 1940 : data_o = 23'b 11010111100010110000100 ;
		12'd 1941 : data_o = 23'b 11010111011000110000101 ;
		12'd 1942 : data_o = 23'b 11010111001110110001001 ;
		12'd 1943 : data_o = 23'b 11010111000100110010000 ;
		12'd 1944 : data_o = 23'b 11010110111010110011001 ;
		12'd 1945 : data_o = 23'b 11010110110000110100100 ;
		12'd 1946 : data_o = 23'b 11010110100110110110011 ;
		12'd 1947 : data_o = 23'b 11010110011100111000011 ;
		12'd 1948 : data_o = 23'b 11010110010010111010111 ;
		12'd 1949 : data_o = 23'b 11010110001000111101100 ;
		12'd 1950 : data_o = 23'b 11010101111111000000101 ;
		12'd 1951 : data_o = 23'b 11010101110101000100000 ;
		12'd 1952 : data_o = 23'b 11010101101011000111101 ;
		12'd 1953 : data_o = 23'b 11010101100001001011101 ;
		12'd 1954 : data_o = 23'b 11010101010111001111111 ;
		12'd 1955 : data_o = 23'b 11010101001101010100100 ;
		12'd 1956 : data_o = 23'b 11010101000011011001100 ;
		12'd 1957 : data_o = 23'b 11010100111001011110110 ;
		12'd 1958 : data_o = 23'b 11010100101111100100010 ;
		12'd 1959 : data_o = 23'b 11010100100101101010001 ;
		12'd 1960 : data_o = 23'b 11010100011011110000011 ;
		12'd 1961 : data_o = 23'b 11010100010001110110111 ;
		12'd 1962 : data_o = 23'b 11010100000111111101101 ;
		12'd 1963 : data_o = 23'b 11010011111110000100110 ;
		12'd 1964 : data_o = 23'b 11010011110100001100010 ;
		12'd 1965 : data_o = 23'b 11010011101010010100000 ;
		12'd 1966 : data_o = 23'b 11010011100000011100000 ;
		12'd 1967 : data_o = 23'b 11010011010110100100011 ;
		12'd 1968 : data_o = 23'b 11010011001100101101001 ;
		12'd 1969 : data_o = 23'b 11010011000010110110001 ;
		12'd 1970 : data_o = 23'b 11010010111000111111100 ;
		12'd 1971 : data_o = 23'b 11010010101111001001001 ;
		12'd 1972 : data_o = 23'b 11010010100101010011000 ;
		12'd 1973 : data_o = 23'b 11010010011011011101010 ;
		12'd 1974 : data_o = 23'b 11010010010001100111111 ;
		12'd 1975 : data_o = 23'b 11010010000111110010110 ;
		12'd 1976 : data_o = 23'b 11010001111101111101111 ;
		12'd 1977 : data_o = 23'b 11010001110100001001011 ;
		12'd 1978 : data_o = 23'b 11010001101010010101010 ;
		12'd 1979 : data_o = 23'b 11010001100000100001011 ;
		12'd 1980 : data_o = 23'b 11010001010110101101110 ;
		12'd 1981 : data_o = 23'b 11010001001100111010100 ;
		12'd 1982 : data_o = 23'b 11010001000011000111100 ;
		12'd 1983 : data_o = 23'b 11010000111001010100111 ;
		12'd 1984 : data_o = 23'b 11010000101111100010100 ;
		12'd 1985 : data_o = 23'b 11010000100101110000100 ;
		12'd 1986 : data_o = 23'b 11010000011011111110110 ;
		12'd 1987 : data_o = 23'b 11010000010010001101011 ;
		12'd 1988 : data_o = 23'b 11010000001000011100010 ;
		12'd 1989 : data_o = 23'b 11001111111110101011100 ;
		12'd 1990 : data_o = 23'b 11001111110100111011000 ;
		12'd 1991 : data_o = 23'b 11001111101011001010111 ;
		12'd 1992 : data_o = 23'b 11001111100001011011000 ;
		12'd 1993 : data_o = 23'b 11001111010111101011011 ;
		12'd 1994 : data_o = 23'b 11001111001101111100001 ;
		12'd 1995 : data_o = 23'b 11001111000100001101010 ;
		12'd 1996 : data_o = 23'b 11001110111010011110101 ;
		12'd 1997 : data_o = 23'b 11001110110000110000010 ;
		12'd 1998 : data_o = 23'b 11001110100111000010010 ;
		12'd 1999 : data_o = 23'b 11001110011101010100100 ;
		12'd 2000 : data_o = 23'b 11001110010011100111001 ;
		12'd 2001 : data_o = 23'b 11001110001001111010000 ;
		12'd 2002 : data_o = 23'b 11001110000000001101001 ;
		12'd 2003 : data_o = 23'b 11001101110110100000101 ;
		12'd 2004 : data_o = 23'b 11001101101100110100100 ;
		12'd 2005 : data_o = 23'b 11001101100011001000101 ;
		12'd 2006 : data_o = 23'b 11001101011001011101000 ;
		12'd 2007 : data_o = 23'b 11001101001111110001110 ;
		12'd 2008 : data_o = 23'b 11001101000110000110110 ;
		12'd 2009 : data_o = 23'b 11001100111100011100001 ;
		12'd 2010 : data_o = 23'b 11001100110010110001110 ;
		12'd 2011 : data_o = 23'b 11001100101001000111101 ;
		12'd 2012 : data_o = 23'b 11001100011111011101111 ;
		12'd 2013 : data_o = 23'b 11001100010101110100011 ;
		12'd 2014 : data_o = 23'b 11001100001100001011010 ;
		12'd 2015 : data_o = 23'b 11001100000010100010011 ;
		12'd 2016 : data_o = 23'b 11001011111000111001111 ;
		12'd 2017 : data_o = 23'b 11001011101111010001101 ;
		12'd 2018 : data_o = 23'b 11001011100101101001110 ;
		12'd 2019 : data_o = 23'b 11001011011100000010000 ;
		12'd 2020 : data_o = 23'b 11001011010010011010110 ;
		12'd 2021 : data_o = 23'b 11001011001000110011101 ;
		12'd 2022 : data_o = 23'b 11001010111111001101000 ;
		12'd 2023 : data_o = 23'b 11001010110101100110100 ;
		12'd 2024 : data_o = 23'b 11001010101100000000011 ;
		12'd 2025 : data_o = 23'b 11001010100010011010100 ;
		12'd 2026 : data_o = 23'b 11001010011000110101000 ;
		12'd 2027 : data_o = 23'b 11001010001111001111110 ;
		12'd 2028 : data_o = 23'b 11001010000101101010111 ;
		12'd 2029 : data_o = 23'b 11001001111100000110010 ;
		12'd 2030 : data_o = 23'b 11001001110010100001111 ;
		12'd 2031 : data_o = 23'b 11001001101000111101111 ;
		12'd 2032 : data_o = 23'b 11001001011111011010001 ;
		12'd 2033 : data_o = 23'b 11001001010101110110110 ;
		12'd 2034 : data_o = 23'b 11001001001100010011101 ;
		12'd 2035 : data_o = 23'b 11001001000010110000110 ;
		12'd 2036 : data_o = 23'b 11001000111001001110010 ;
		12'd 2037 : data_o = 23'b 11001000101111101100000 ;
		12'd 2038 : data_o = 23'b 11001000100110001010000 ;
		12'd 2039 : data_o = 23'b 11001000011100101000011 ;
		12'd 2040 : data_o = 23'b 11001000010011000111001 ;
		12'd 2041 : data_o = 23'b 11001000001001100110000 ;
		12'd 2042 : data_o = 23'b 11001000000000000101010 ;
		12'd 2043 : data_o = 23'b 11000111110110100100111 ;
		12'd 2044 : data_o = 23'b 11000111101101000100101 ;
		12'd 2045 : data_o = 23'b 11000111100011100100111 ;
		12'd 2046 : data_o = 23'b 11000111011010000101010 ;
		12'd 2047 : data_o = 23'b 11000111010000100110000 ;
		12'd 2048 : data_o = 23'b 11000111000111000111000 ;
		12'd 2049 : data_o = 23'b 11000110111101101000011 ;
		12'd 2050 : data_o = 23'b 11000110110100001010000 ;
		12'd 2051 : data_o = 23'b 11000110101010101011111 ;
		12'd 2052 : data_o = 23'b 11000110100001001110001 ;
		12'd 2053 : data_o = 23'b 11000110010111110000101 ;
		12'd 2054 : data_o = 23'b 11000110001110010011100 ;
		12'd 2055 : data_o = 23'b 11000110000100110110101 ;
		12'd 2056 : data_o = 23'b 11000101111011011010000 ;
		12'd 2057 : data_o = 23'b 11000101110001111101110 ;
		12'd 2058 : data_o = 23'b 11000101101000100001101 ;
		12'd 2059 : data_o = 23'b 11000101011111000110000 ;
		12'd 2060 : data_o = 23'b 11000101010101101010100 ;
		12'd 2061 : data_o = 23'b 11000101001100001111011 ;
		12'd 2062 : data_o = 23'b 11000101000010110100101 ;
		12'd 2063 : data_o = 23'b 11000100111001011010000 ;
		12'd 2064 : data_o = 23'b 11000100101111111111110 ;
		12'd 2065 : data_o = 23'b 11000100100110100101111 ;
		12'd 2066 : data_o = 23'b 11000100011101001100010 ;
		12'd 2067 : data_o = 23'b 11000100010011110010111 ;
		12'd 2068 : data_o = 23'b 11000100001010011001110 ;
		12'd 2069 : data_o = 23'b 11000100000001000001000 ;
		12'd 2070 : data_o = 23'b 11000011110111101000100 ;
		12'd 2071 : data_o = 23'b 11000011101110010000010 ;
		12'd 2072 : data_o = 23'b 11000011100100111000011 ;
		12'd 2073 : data_o = 23'b 11000011011011100000110 ;
		12'd 2074 : data_o = 23'b 11000011010010001001100 ;
		12'd 2075 : data_o = 23'b 11000011001000110010011 ;
		12'd 2076 : data_o = 23'b 11000010111111011011101 ;
		12'd 2077 : data_o = 23'b 11000010110110000101010 ;
		12'd 2078 : data_o = 23'b 11000010101100101111001 ;
		12'd 2079 : data_o = 23'b 11000010100011011001010 ;
		12'd 2080 : data_o = 23'b 11000010011010000011101 ;
		12'd 2081 : data_o = 23'b 11000010010000101110011 ;
		12'd 2082 : data_o = 23'b 11000010000111011001011 ;
		12'd 2083 : data_o = 23'b 11000001111110000100101 ;
		12'd 2084 : data_o = 23'b 11000001110100110000010 ;
		12'd 2085 : data_o = 23'b 11000001101011011100001 ;
		12'd 2086 : data_o = 23'b 11000001100010001000010 ;
		12'd 2087 : data_o = 23'b 11000001011000110100110 ;
		12'd 2088 : data_o = 23'b 11000001001111100001100 ;
		12'd 2089 : data_o = 23'b 11000001000110001110100 ;
		12'd 2090 : data_o = 23'b 11000000111100111011110 ;
		12'd 2091 : data_o = 23'b 11000000110011101001011 ;
		12'd 2092 : data_o = 23'b 11000000101010010111010 ;
		12'd 2093 : data_o = 23'b 11000000100001000101100 ;
		12'd 2094 : data_o = 23'b 11000000010111110100000 ;
		12'd 2095 : data_o = 23'b 11000000001110100010110 ;
		12'd 2096 : data_o = 23'b 11000000000101010001110 ;
		12'd 2097 : data_o = 23'b 10111111111100000001001 ;
		12'd 2098 : data_o = 23'b 10111111110010110000110 ;
		12'd 2099 : data_o = 23'b 10111111101001100000101 ;
		12'd 2100 : data_o = 23'b 10111111100000010000110 ;
		12'd 2101 : data_o = 23'b 10111111010111000001010 ;
		12'd 2102 : data_o = 23'b 10111111001101110010000 ;
		12'd 2103 : data_o = 23'b 10111111000100100011001 ;
		12'd 2104 : data_o = 23'b 10111110111011010100011 ;
		12'd 2105 : data_o = 23'b 10111110110010000110000 ;
		12'd 2106 : data_o = 23'b 10111110101000111000000 ;
		12'd 2107 : data_o = 23'b 10111110011111101010001 ;
		12'd 2108 : data_o = 23'b 10111110010110011100101 ;
		12'd 2109 : data_o = 23'b 10111110001101001111011 ;
		12'd 2110 : data_o = 23'b 10111110000100000010100 ;
		12'd 2111 : data_o = 23'b 10111101111010110101110 ;
		12'd 2112 : data_o = 23'b 10111101110001101001011 ;
		12'd 2113 : data_o = 23'b 10111101101000011101010 ;
		12'd 2114 : data_o = 23'b 10111101011111010001100 ;
		12'd 2115 : data_o = 23'b 10111101010110000110000 ;
		12'd 2116 : data_o = 23'b 10111101001100111010110 ;
		12'd 2117 : data_o = 23'b 10111101000011101111110 ;
		12'd 2118 : data_o = 23'b 10111100111010100101001 ;
		12'd 2119 : data_o = 23'b 10111100110001011010101 ;
		12'd 2120 : data_o = 23'b 10111100101000010000100 ;
		12'd 2121 : data_o = 23'b 10111100011111000110110 ;
		12'd 2122 : data_o = 23'b 10111100010101111101001 ;
		12'd 2123 : data_o = 23'b 10111100001100110011111 ;
		12'd 2124 : data_o = 23'b 10111100000011101010111 ;
		12'd 2125 : data_o = 23'b 10111011111010100010010 ;
		12'd 2126 : data_o = 23'b 10111011110001011001110 ;
		12'd 2127 : data_o = 23'b 10111011101000010001101 ;
		12'd 2128 : data_o = 23'b 10111011011111001001111 ;
		12'd 2129 : data_o = 23'b 10111011010110000010010 ;
		12'd 2130 : data_o = 23'b 10111011001100111011000 ;
		12'd 2131 : data_o = 23'b 10111011000011110011111 ;
		12'd 2132 : data_o = 23'b 10111010111010101101010 ;
		12'd 2133 : data_o = 23'b 10111010110001100110110 ;
		12'd 2134 : data_o = 23'b 10111010101000100000101 ;
		12'd 2135 : data_o = 23'b 10111010011111011010110 ;
		12'd 2136 : data_o = 23'b 10111010010110010101001 ;
		12'd 2137 : data_o = 23'b 10111010001101001111110 ;
		12'd 2138 : data_o = 23'b 10111010000100001010110 ;
		12'd 2139 : data_o = 23'b 10111001111011000101111 ;
		12'd 2140 : data_o = 23'b 10111001110010000001011 ;
		12'd 2141 : data_o = 23'b 10111001101000111101010 ;
		12'd 2142 : data_o = 23'b 10111001011111111001010 ;
		12'd 2143 : data_o = 23'b 10111001010110110101101 ;
		12'd 2144 : data_o = 23'b 10111001001101110010010 ;
		12'd 2145 : data_o = 23'b 10111001000100101111001 ;
		12'd 2146 : data_o = 23'b 10111000111011101100011 ;
		12'd 2147 : data_o = 23'b 10111000110010101001110 ;
		12'd 2148 : data_o = 23'b 10111000101001100111100 ;
		12'd 2149 : data_o = 23'b 10111000100000100101100 ;
		12'd 2150 : data_o = 23'b 10111000010111100011111 ;
		12'd 2151 : data_o = 23'b 10111000001110100010011 ;
		12'd 2152 : data_o = 23'b 10111000000101100001010 ;
		12'd 2153 : data_o = 23'b 10110111111100100000011 ;
		12'd 2154 : data_o = 23'b 10110111110011011111110 ;
		12'd 2155 : data_o = 23'b 10110111101010011111100 ;
		12'd 2156 : data_o = 23'b 10110111100001011111011 ;
		12'd 2157 : data_o = 23'b 10110111011000011111101 ;
		12'd 2158 : data_o = 23'b 10110111001111100000001 ;
		12'd 2159 : data_o = 23'b 10110111000110100001000 ;
		12'd 2160 : data_o = 23'b 10110110111101100010000 ;
		12'd 2161 : data_o = 23'b 10110110110100100011011 ;
		12'd 2162 : data_o = 23'b 10110110101011100101000 ;
		12'd 2163 : data_o = 23'b 10110110100010100110111 ;
		12'd 2164 : data_o = 23'b 10110110011001101001000 ;
		12'd 2165 : data_o = 23'b 10110110010000101011011 ;
		12'd 2166 : data_o = 23'b 10110110000111101110001 ;
		12'd 2167 : data_o = 23'b 10110101111110110001001 ;
		12'd 2168 : data_o = 23'b 10110101110101110100011 ;
		12'd 2169 : data_o = 23'b 10110101101100110111111 ;
		12'd 2170 : data_o = 23'b 10110101100011111011110 ;
		12'd 2171 : data_o = 23'b 10110101011010111111110 ;
		12'd 2172 : data_o = 23'b 10110101010010000100001 ;
		12'd 2173 : data_o = 23'b 10110101001001001000110 ;
		12'd 2174 : data_o = 23'b 10110101000000001101101 ;
		12'd 2175 : data_o = 23'b 10110100110111010010111 ;
		12'd 2176 : data_o = 23'b 10110100101110011000010 ;
		12'd 2177 : data_o = 23'b 10110100100101011110000 ;
		12'd 2178 : data_o = 23'b 10110100011100100100000 ;
		12'd 2179 : data_o = 23'b 10110100010011101010010 ;
		12'd 2180 : data_o = 23'b 10110100001010110000111 ;
		12'd 2181 : data_o = 23'b 10110100000001110111101 ;
		12'd 2182 : data_o = 23'b 10110011111000111110110 ;
		12'd 2183 : data_o = 23'b 10110011110000000110001 ;
		12'd 2184 : data_o = 23'b 10110011100111001101110 ;
		12'd 2185 : data_o = 23'b 10110011011110010101101 ;
		12'd 2186 : data_o = 23'b 10110011010101011101110 ;
		12'd 2187 : data_o = 23'b 10110011001100100110010 ;
		12'd 2188 : data_o = 23'b 10110011000011101110111 ;
		12'd 2189 : data_o = 23'b 10110010111010110111111 ;
		12'd 2190 : data_o = 23'b 10110010110010000001001 ;
		12'd 2191 : data_o = 23'b 10110010101001001010101 ;
		12'd 2192 : data_o = 23'b 10110010100000010100100 ;
		12'd 2193 : data_o = 23'b 10110010010111011110100 ;
		12'd 2194 : data_o = 23'b 10110010001110101000111 ;
		12'd 2195 : data_o = 23'b 10110010000101110011100 ;
		12'd 2196 : data_o = 23'b 10110001111100111110011 ;
		12'd 2197 : data_o = 23'b 10110001110100001001100 ;
		12'd 2198 : data_o = 23'b 10110001101011010100111 ;
		12'd 2199 : data_o = 23'b 10110001100010100000100 ;
		12'd 2200 : data_o = 23'b 10110001011001101100100 ;
		12'd 2201 : data_o = 23'b 10110001010000111000110 ;
		12'd 2202 : data_o = 23'b 10110001001000000101010 ;
		12'd 2203 : data_o = 23'b 10110000111111010010000 ;
		12'd 2204 : data_o = 23'b 10110000110110011111000 ;
		12'd 2205 : data_o = 23'b 10110000101101101100010 ;
		12'd 2206 : data_o = 23'b 10110000100100111001111 ;
		12'd 2207 : data_o = 23'b 10110000011100000111101 ;
		12'd 2208 : data_o = 23'b 10110000010011010101110 ;
		12'd 2209 : data_o = 23'b 10110000001010100100001 ;
		12'd 2210 : data_o = 23'b 10110000000001110010110 ;
		12'd 2211 : data_o = 23'b 10101111111001000001101 ;
		12'd 2212 : data_o = 23'b 10101111110000010000110 ;
		12'd 2213 : data_o = 23'b 10101111100111100000010 ;
		12'd 2214 : data_o = 23'b 10101111011110101111111 ;
		12'd 2215 : data_o = 23'b 10101111010101111111111 ;
		12'd 2216 : data_o = 23'b 10101111001101010000001 ;
		12'd 2217 : data_o = 23'b 10101111000100100000101 ;
		12'd 2218 : data_o = 23'b 10101110111011110001011 ;
		12'd 2219 : data_o = 23'b 10101110110011000010011 ;
		12'd 2220 : data_o = 23'b 10101110101010010011101 ;
		12'd 2221 : data_o = 23'b 10101110100001100101010 ;
		12'd 2222 : data_o = 23'b 10101110011000110111000 ;
		12'd 2223 : data_o = 23'b 10101110010000001001001 ;
		12'd 2224 : data_o = 23'b 10101110000111011011100 ;
		12'd 2225 : data_o = 23'b 10101101111110101110001 ;
		12'd 2226 : data_o = 23'b 10101101110110000001000 ;
		12'd 2227 : data_o = 23'b 10101101101101010100001 ;
		12'd 2228 : data_o = 23'b 10101101100100100111100 ;
		12'd 2229 : data_o = 23'b 10101101011011111011001 ;
		12'd 2230 : data_o = 23'b 10101101010011001111001 ;
		12'd 2231 : data_o = 23'b 10101101001010100011011 ;
		12'd 2232 : data_o = 23'b 10101101000001110111110 ;
		12'd 2233 : data_o = 23'b 10101100111001001100100 ;
		12'd 2234 : data_o = 23'b 10101100110000100001100 ;
		12'd 2235 : data_o = 23'b 10101100100111110110110 ;
		12'd 2236 : data_o = 23'b 10101100011111001100010 ;
		12'd 2237 : data_o = 23'b 10101100010110100010000 ;
		12'd 2238 : data_o = 23'b 10101100001101111000001 ;
		12'd 2239 : data_o = 23'b 10101100000101001110011 ;
		12'd 2240 : data_o = 23'b 10101011111100100101000 ;
		12'd 2241 : data_o = 23'b 10101011110011111011110 ;
		12'd 2242 : data_o = 23'b 10101011101011010010111 ;
		12'd 2243 : data_o = 23'b 10101011100010101010010 ;
		12'd 2244 : data_o = 23'b 10101011011010000001111 ;
		12'd 2245 : data_o = 23'b 10101011010001011001110 ;
		12'd 2246 : data_o = 23'b 10101011001000110001111 ;
		12'd 2247 : data_o = 23'b 10101011000000001010010 ;
		12'd 2248 : data_o = 23'b 10101010110111100010111 ;
		12'd 2249 : data_o = 23'b 10101010101110111011110 ;
		12'd 2250 : data_o = 23'b 10101010100110010101000 ;
		12'd 2251 : data_o = 23'b 10101010011101101110011 ;
		12'd 2252 : data_o = 23'b 10101010010101001000001 ;
		12'd 2253 : data_o = 23'b 10101010001100100010001 ;
		12'd 2254 : data_o = 23'b 10101010000011111100010 ;
		12'd 2255 : data_o = 23'b 10101001111011010110110 ;
		12'd 2256 : data_o = 23'b 10101001110010110001100 ;
		12'd 2257 : data_o = 23'b 10101001101010001100100 ;
		12'd 2258 : data_o = 23'b 10101001100001100111110 ;
		12'd 2259 : data_o = 23'b 10101001011001000011010 ;
		12'd 2260 : data_o = 23'b 10101001010000011111000 ;
		12'd 2261 : data_o = 23'b 10101001000111111011001 ;
		12'd 2262 : data_o = 23'b 10101000111111010111011 ;
		12'd 2263 : data_o = 23'b 10101000110110110011111 ;
		12'd 2264 : data_o = 23'b 10101000101110010000110 ;
		12'd 2265 : data_o = 23'b 10101000100101101101110 ;
		12'd 2266 : data_o = 23'b 10101000011101001011001 ;
		12'd 2267 : data_o = 23'b 10101000010100101000101 ;
		12'd 2268 : data_o = 23'b 10101000001100000110100 ;
		12'd 2269 : data_o = 23'b 10101000000011100100101 ;
		12'd 2270 : data_o = 23'b 10100111111011000011000 ;
		12'd 2271 : data_o = 23'b 10100111110010100001101 ;
		12'd 2272 : data_o = 23'b 10100111101010000000100 ;
		12'd 2273 : data_o = 23'b 10100111100001011111100 ;
		12'd 2274 : data_o = 23'b 10100111011000111111000 ;
		12'd 2275 : data_o = 23'b 10100111010000011110101 ;
		12'd 2276 : data_o = 23'b 10100111000111111110100 ;
		12'd 2277 : data_o = 23'b 10100110111111011110101 ;
		12'd 2278 : data_o = 23'b 10100110110110111111000 ;
		12'd 2279 : data_o = 23'b 10100110101110011111101 ;
		12'd 2280 : data_o = 23'b 10100110100110000000101 ;
		12'd 2281 : data_o = 23'b 10100110011101100001110 ;
		12'd 2282 : data_o = 23'b 10100110010101000011010 ;
		12'd 2283 : data_o = 23'b 10100110001100100100111 ;
		12'd 2284 : data_o = 23'b 10100110000100000110111 ;
		12'd 2285 : data_o = 23'b 10100101111011101001000 ;
		12'd 2286 : data_o = 23'b 10100101110011001011100 ;
		12'd 2287 : data_o = 23'b 10100101101010101110001 ;
		12'd 2288 : data_o = 23'b 10100101100010010001001 ;
		12'd 2289 : data_o = 23'b 10100101011001110100011 ;
		12'd 2290 : data_o = 23'b 10100101010001010111110 ;
		12'd 2291 : data_o = 23'b 10100101001000111011100 ;
		12'd 2292 : data_o = 23'b 10100101000000011111100 ;
		12'd 2293 : data_o = 23'b 10100100111000000011110 ;
		12'd 2294 : data_o = 23'b 10100100101111101000001 ;
		12'd 2295 : data_o = 23'b 10100100100111001100111 ;
		12'd 2296 : data_o = 23'b 10100100011110110001111 ;
		12'd 2297 : data_o = 23'b 10100100010110010111001 ;
		12'd 2298 : data_o = 23'b 10100100001101111100101 ;
		12'd 2299 : data_o = 23'b 10100100000101100010011 ;
		12'd 2300 : data_o = 23'b 10100011111101001000011 ;
		12'd 2301 : data_o = 23'b 10100011110100101110101 ;
		12'd 2302 : data_o = 23'b 10100011101100010101001 ;
		12'd 2303 : data_o = 23'b 10100011100011111011111 ;
		12'd 2304 : data_o = 23'b 10100011011011100010111 ;
		12'd 2305 : data_o = 23'b 10100011010011001010001 ;
		12'd 2306 : data_o = 23'b 10100011001010110001101 ;
		12'd 2307 : data_o = 23'b 10100011000010011001011 ;
		12'd 2308 : data_o = 23'b 10100010111010000001011 ;
		12'd 2309 : data_o = 23'b 10100010110001101001101 ;
		12'd 2310 : data_o = 23'b 10100010101001010010001 ;
		12'd 2311 : data_o = 23'b 10100010100000111010111 ;
		12'd 2312 : data_o = 23'b 10100010011000100011111 ;
		12'd 2313 : data_o = 23'b 10100010010000001101010 ;
		12'd 2314 : data_o = 23'b 10100010000111110110110 ;
		12'd 2315 : data_o = 23'b 10100001111111100000100 ;
		12'd 2316 : data_o = 23'b 10100001110111001010100 ;
		12'd 2317 : data_o = 23'b 10100001101110110100110 ;
		12'd 2318 : data_o = 23'b 10100001100110011111010 ;
		12'd 2319 : data_o = 23'b 10100001011110001010000 ;
		12'd 2320 : data_o = 23'b 10100001010101110101000 ;
		12'd 2321 : data_o = 23'b 10100001001101100000010 ;
		12'd 2322 : data_o = 23'b 10100001000101001011110 ;
		12'd 2323 : data_o = 23'b 10100000111100110111100 ;
		12'd 2324 : data_o = 23'b 10100000110100100011100 ;
		12'd 2325 : data_o = 23'b 10100000101100001111111 ;
		12'd 2326 : data_o = 23'b 10100000100011111100011 ;
		12'd 2327 : data_o = 23'b 10100000011011101001001 ;
		12'd 2328 : data_o = 23'b 10100000010011010110001 ;
		12'd 2329 : data_o = 23'b 10100000001011000011011 ;
		12'd 2330 : data_o = 23'b 10100000000010110000111 ;
		12'd 2331 : data_o = 23'b 10011111111010011110100 ;
		12'd 2332 : data_o = 23'b 10011111110010001100100 ;
		12'd 2333 : data_o = 23'b 10011111101001111010110 ;
		12'd 2334 : data_o = 23'b 10011111100001101001010 ;
		12'd 2335 : data_o = 23'b 10011111011001011000000 ;
		12'd 2336 : data_o = 23'b 10011111010001000111000 ;
		12'd 2337 : data_o = 23'b 10011111001000110110010 ;
		12'd 2338 : data_o = 23'b 10011111000000100101101 ;
		12'd 2339 : data_o = 23'b 10011110111000010101011 ;
		12'd 2340 : data_o = 23'b 10011110110000000101011 ;
		12'd 2341 : data_o = 23'b 10011110100111110101101 ;
		12'd 2342 : data_o = 23'b 10011110011111100110000 ;
		12'd 2343 : data_o = 23'b 10011110010111010110110 ;
		12'd 2344 : data_o = 23'b 10011110001111000111101 ;
		12'd 2345 : data_o = 23'b 10011110000110111000111 ;
		12'd 2346 : data_o = 23'b 10011101111110101010011 ;
		12'd 2347 : data_o = 23'b 10011101110110011100000 ;
		12'd 2348 : data_o = 23'b 10011101101110001101111 ;
		12'd 2349 : data_o = 23'b 10011101100110000000001 ;
		12'd 2350 : data_o = 23'b 10011101011101110010100 ;
		12'd 2351 : data_o = 23'b 10011101010101100101001 ;
		12'd 2352 : data_o = 23'b 10011101001101011000001 ;
		12'd 2353 : data_o = 23'b 10011101000101001011010 ;
		12'd 2354 : data_o = 23'b 10011100111100111110101 ;
		12'd 2355 : data_o = 23'b 10011100110100110010010 ;
		12'd 2356 : data_o = 23'b 10011100101100100110001 ;
		12'd 2357 : data_o = 23'b 10011100100100011010010 ;
		12'd 2358 : data_o = 23'b 10011100011100001110101 ;
		12'd 2359 : data_o = 23'b 10011100010100000011010 ;
		12'd 2360 : data_o = 23'b 10011100001011111000001 ;
		12'd 2361 : data_o = 23'b 10011100000011101101010 ;
		12'd 2362 : data_o = 23'b 10011011111011100010101 ;
		12'd 2363 : data_o = 23'b 10011011110011011000001 ;
		12'd 2364 : data_o = 23'b 10011011101011001110000 ;
		12'd 2365 : data_o = 23'b 10011011100011000100000 ;
		12'd 2366 : data_o = 23'b 10011011011010111010011 ;
		12'd 2367 : data_o = 23'b 10011011010010110000111 ;
		12'd 2368 : data_o = 23'b 10011011001010100111110 ;
		12'd 2369 : data_o = 23'b 10011011000010011110110 ;
		12'd 2370 : data_o = 23'b 10011010111010010110000 ;
		12'd 2371 : data_o = 23'b 10011010110010001101101 ;
		12'd 2372 : data_o = 23'b 10011010101010000101011 ;
		12'd 2373 : data_o = 23'b 10011010100001111101011 ;
		12'd 2374 : data_o = 23'b 10011010011001110101101 ;
		12'd 2375 : data_o = 23'b 10011010010001101110001 ;
		12'd 2376 : data_o = 23'b 10011010001001100110110 ;
		12'd 2377 : data_o = 23'b 10011010000001011111110 ;
		12'd 2378 : data_o = 23'b 10011001111001011001000 ;
		12'd 2379 : data_o = 23'b 10011001110001010010011 ;
		12'd 2380 : data_o = 23'b 10011001101001001100001 ;
		12'd 2381 : data_o = 23'b 10011001100001000110000 ;
		12'd 2382 : data_o = 23'b 10011001011001000000010 ;
		12'd 2383 : data_o = 23'b 10011001010000111010101 ;
		12'd 2384 : data_o = 23'b 10011001001000110101010 ;
		12'd 2385 : data_o = 23'b 10011001000000110000001 ;
		12'd 2386 : data_o = 23'b 10011000111000101011010 ;
		12'd 2387 : data_o = 23'b 10011000110000100110101 ;
		12'd 2388 : data_o = 23'b 10011000101000100010010 ;
		12'd 2389 : data_o = 23'b 10011000100000011110001 ;
		12'd 2390 : data_o = 23'b 10011000011000011010010 ;
		12'd 2391 : data_o = 23'b 10011000010000010110100 ;
		12'd 2392 : data_o = 23'b 10011000001000010011001 ;
		12'd 2393 : data_o = 23'b 10011000000000001111111 ;
		12'd 2394 : data_o = 23'b 10010111111000001100111 ;
		12'd 2395 : data_o = 23'b 10010111110000001010001 ;
		12'd 2396 : data_o = 23'b 10010111101000000111110 ;
		12'd 2397 : data_o = 23'b 10010111100000000101100 ;
		12'd 2398 : data_o = 23'b 10010111011000000011011 ;
		12'd 2399 : data_o = 23'b 10010111010000000001101 ;
		12'd 2400 : data_o = 23'b 10010111001000000000001 ;
		12'd 2401 : data_o = 23'b 10010110111111111110111 ;
		12'd 2402 : data_o = 23'b 10010110110111111101110 ;
		12'd 2403 : data_o = 23'b 10010110101111111100111 ;
		12'd 2404 : data_o = 23'b 10010110100111111100011 ;
		12'd 2405 : data_o = 23'b 10010110011111111100000 ;
		12'd 2406 : data_o = 23'b 10010110010111111011111 ;
		12'd 2407 : data_o = 23'b 10010110001111111100000 ;
		12'd 2408 : data_o = 23'b 10010110000111111100011 ;
		12'd 2409 : data_o = 23'b 10010101111111111101000 ;
		12'd 2410 : data_o = 23'b 10010101110111111101110 ;
		12'd 2411 : data_o = 23'b 10010101101111111110111 ;
		12'd 2412 : data_o = 23'b 10010101101000000000001 ;
		12'd 2413 : data_o = 23'b 10010101100000000001101 ;
		12'd 2414 : data_o = 23'b 10010101011000000011011 ;
		12'd 2415 : data_o = 23'b 10010101010000000101011 ;
		12'd 2416 : data_o = 23'b 10010101001000000111101 ;
		12'd 2417 : data_o = 23'b 10010101000000001010001 ;
		12'd 2418 : data_o = 23'b 10010100111000001100111 ;
		12'd 2419 : data_o = 23'b 10010100110000001111110 ;
		12'd 2420 : data_o = 23'b 10010100101000010011000 ;
		12'd 2421 : data_o = 23'b 10010100100000010110011 ;
		12'd 2422 : data_o = 23'b 10010100011000011010000 ;
		12'd 2423 : data_o = 23'b 10010100010000011101111 ;
		12'd 2424 : data_o = 23'b 10010100001000100010000 ;
		12'd 2425 : data_o = 23'b 10010100000000100110011 ;
		12'd 2426 : data_o = 23'b 10010011111000101011000 ;
		12'd 2427 : data_o = 23'b 10010011110000101111110 ;
		12'd 2428 : data_o = 23'b 10010011101000110100111 ;
		12'd 2429 : data_o = 23'b 10010011100000111010001 ;
		12'd 2430 : data_o = 23'b 10010011011000111111101 ;
		12'd 2431 : data_o = 23'b 10010011010001000101011 ;
		12'd 2432 : data_o = 23'b 10010011001001001011011 ;
		12'd 2433 : data_o = 23'b 10010011000001010001100 ;
		12'd 2434 : data_o = 23'b 10010010111001011000000 ;
		12'd 2435 : data_o = 23'b 10010010110001011110101 ;
		12'd 2436 : data_o = 23'b 10010010101001100101101 ;
		12'd 2437 : data_o = 23'b 10010010100001101100110 ;
		12'd 2438 : data_o = 23'b 10010010011001110100001 ;
		12'd 2439 : data_o = 23'b 10010010010001111011101 ;
		12'd 2440 : data_o = 23'b 10010010001010000011100 ;
		12'd 2441 : data_o = 23'b 10010010000010001011101 ;
		12'd 2442 : data_o = 23'b 10010001111010010011111 ;
		12'd 2443 : data_o = 23'b 10010001110010011100011 ;
		12'd 2444 : data_o = 23'b 10010001101010100101001 ;
		12'd 2445 : data_o = 23'b 10010001100010101110001 ;
		12'd 2446 : data_o = 23'b 10010001011010110111011 ;
		12'd 2447 : data_o = 23'b 10010001010011000000111 ;
		12'd 2448 : data_o = 23'b 10010001001011001010100 ;
		12'd 2449 : data_o = 23'b 10010001000011010100011 ;
		12'd 2450 : data_o = 23'b 10010000111011011110100 ;
		12'd 2451 : data_o = 23'b 10010000110011101000111 ;
		12'd 2452 : data_o = 23'b 10010000101011110011100 ;
		12'd 2453 : data_o = 23'b 10010000100011111110011 ;
		12'd 2454 : data_o = 23'b 10010000011100001001011 ;
		12'd 2455 : data_o = 23'b 10010000010100010100110 ;
		12'd 2456 : data_o = 23'b 10010000001100100000010 ;
		12'd 2457 : data_o = 23'b 10010000000100101100000 ;
		12'd 2458 : data_o = 23'b 10001111111100111000000 ;
		12'd 2459 : data_o = 23'b 10001111110101000100001 ;
		12'd 2460 : data_o = 23'b 10001111101101010000101 ;
		12'd 2461 : data_o = 23'b 10001111100101011101010 ;
		12'd 2462 : data_o = 23'b 10001111011101101010001 ;
		12'd 2463 : data_o = 23'b 10001111010101110111010 ;
		12'd 2464 : data_o = 23'b 10001111001110000100101 ;
		12'd 2465 : data_o = 23'b 10001111000110010010010 ;
		12'd 2466 : data_o = 23'b 10001110111110100000000 ;
		12'd 2467 : data_o = 23'b 10001110110110101110000 ;
		12'd 2468 : data_o = 23'b 10001110101110111100010 ;
		12'd 2469 : data_o = 23'b 10001110100111001010110 ;
		12'd 2470 : data_o = 23'b 10001110011111011001100 ;
		12'd 2471 : data_o = 23'b 10001110010111101000011 ;
		12'd 2472 : data_o = 23'b 10001110001111110111101 ;
		12'd 2473 : data_o = 23'b 10001110001000000111000 ;
		12'd 2474 : data_o = 23'b 10001110000000010110101 ;
		12'd 2475 : data_o = 23'b 10001101111000100110100 ;
		12'd 2476 : data_o = 23'b 10001101110000110110100 ;
		12'd 2477 : data_o = 23'b 10001101101001000110111 ;
		12'd 2478 : data_o = 23'b 10001101100001010111011 ;
		12'd 2479 : data_o = 23'b 10001101011001101000001 ;
		12'd 2480 : data_o = 23'b 10001101010001111001001 ;
		12'd 2481 : data_o = 23'b 10001101001010001010010 ;
		12'd 2482 : data_o = 23'b 10001101000010011011110 ;
		12'd 2483 : data_o = 23'b 10001100111010101101011 ;
		12'd 2484 : data_o = 23'b 10001100110010111111010 ;
		12'd 2485 : data_o = 23'b 10001100101011010001011 ;
		12'd 2486 : data_o = 23'b 10001100100011100011110 ;
		12'd 2487 : data_o = 23'b 10001100011011110110010 ;
		12'd 2488 : data_o = 23'b 10001100010100001001000 ;
		12'd 2489 : data_o = 23'b 10001100001100011100000 ;
		12'd 2490 : data_o = 23'b 10001100000100101111010 ;
		12'd 2491 : data_o = 23'b 10001011111101000010110 ;
		12'd 2492 : data_o = 23'b 10001011110101010110011 ;
		12'd 2493 : data_o = 23'b 10001011101101101010011 ;
		12'd 2494 : data_o = 23'b 10001011100101111110100 ;
		12'd 2495 : data_o = 23'b 10001011011110010010110 ;
		12'd 2496 : data_o = 23'b 10001011010110100111011 ;
		12'd 2497 : data_o = 23'b 10001011001110111100001 ;
		12'd 2498 : data_o = 23'b 10001011000111010001010 ;
		12'd 2499 : data_o = 23'b 10001010111111100110100 ;
		12'd 2500 : data_o = 23'b 10001010110111111011111 ;
		12'd 2501 : data_o = 23'b 10001010110000010001101 ;
		12'd 2502 : data_o = 23'b 10001010101000100111100 ;
		12'd 2503 : data_o = 23'b 10001010100000111101101 ;
		12'd 2504 : data_o = 23'b 10001010011001010100000 ;
		12'd 2505 : data_o = 23'b 10001010010001101010101 ;
		12'd 2506 : data_o = 23'b 10001010001010000001011 ;
		12'd 2507 : data_o = 23'b 10001010000010011000011 ;
		12'd 2508 : data_o = 23'b 10001001111010101111101 ;
		12'd 2509 : data_o = 23'b 10001001110011000111001 ;
		12'd 2510 : data_o = 23'b 10001001101011011110111 ;
		12'd 2511 : data_o = 23'b 10001001100011110110110 ;
		12'd 2512 : data_o = 23'b 10001001011100001110111 ;
		12'd 2513 : data_o = 23'b 10001001010100100111010 ;
		12'd 2514 : data_o = 23'b 10001001001100111111111 ;
		12'd 2515 : data_o = 23'b 10001001000101011000101 ;
		12'd 2516 : data_o = 23'b 10001000111101110001101 ;
		12'd 2517 : data_o = 23'b 10001000110110001010111 ;
		12'd 2518 : data_o = 23'b 10001000101110100100011 ;
		12'd 2519 : data_o = 23'b 10001000100110111110000 ;
		12'd 2520 : data_o = 23'b 10001000011111011000000 ;
		12'd 2521 : data_o = 23'b 10001000010111110010001 ;
		12'd 2522 : data_o = 23'b 10001000010000001100011 ;
		12'd 2523 : data_o = 23'b 10001000001000100111000 ;
		12'd 2524 : data_o = 23'b 10001000000001000001110 ;
		12'd 2525 : data_o = 23'b 10000111111001011100110 ;
		12'd 2526 : data_o = 23'b 10000111110001111000000 ;
		12'd 2527 : data_o = 23'b 10000111101010010011100 ;
		12'd 2528 : data_o = 23'b 10000111100010101111001 ;
		12'd 2529 : data_o = 23'b 10000111011011001011000 ;
		12'd 2530 : data_o = 23'b 10000111010011100111001 ;
		12'd 2531 : data_o = 23'b 10000111001100000011011 ;
		12'd 2532 : data_o = 23'b 10000111000100100000000 ;
		12'd 2533 : data_o = 23'b 10000110111100111100110 ;
		12'd 2534 : data_o = 23'b 10000110110101011001110 ;
		12'd 2535 : data_o = 23'b 10000110101101110110111 ;
		12'd 2536 : data_o = 23'b 10000110100110010100010 ;
		12'd 2537 : data_o = 23'b 10000110011110110001111 ;
		12'd 2538 : data_o = 23'b 10000110010111001111110 ;
		12'd 2539 : data_o = 23'b 10000110001111101101111 ;
		12'd 2540 : data_o = 23'b 10000110001000001100001 ;
		12'd 2541 : data_o = 23'b 10000110000000101010101 ;
		12'd 2542 : data_o = 23'b 10000101111001001001011 ;
		12'd 2543 : data_o = 23'b 10000101110001101000010 ;
		12'd 2544 : data_o = 23'b 10000101101010000111100 ;
		12'd 2545 : data_o = 23'b 10000101100010100110111 ;
		12'd 2546 : data_o = 23'b 10000101011011000110011 ;
		12'd 2547 : data_o = 23'b 10000101010011100110010 ;
		12'd 2548 : data_o = 23'b 10000101001100000110010 ;
		12'd 2549 : data_o = 23'b 10000101000100100110100 ;
		12'd 2550 : data_o = 23'b 10000100111101000111000 ;
		12'd 2551 : data_o = 23'b 10000100110101100111101 ;
		12'd 2552 : data_o = 23'b 10000100101110001000100 ;
		12'd 2553 : data_o = 23'b 10000100100110101001101 ;
		12'd 2554 : data_o = 23'b 10000100011111001011000 ;
		12'd 2555 : data_o = 23'b 10000100010111101100100 ;
		12'd 2556 : data_o = 23'b 10000100010000001110010 ;
		12'd 2557 : data_o = 23'b 10000100001000110000010 ;
		12'd 2558 : data_o = 23'b 10000100000001010010011 ;
		12'd 2559 : data_o = 23'b 10000011111001110100110 ;
		12'd 2560 : data_o = 23'b 10000011110010010111011 ;
		12'd 2561 : data_o = 23'b 10000011101010111010010 ;
		12'd 2562 : data_o = 23'b 10000011100011011101010 ;
		12'd 2563 : data_o = 23'b 10000011011100000000100 ;
		12'd 2564 : data_o = 23'b 10000011010100100100000 ;
		12'd 2565 : data_o = 23'b 10000011001101000111110 ;
		12'd 2566 : data_o = 23'b 10000011000101101011101 ;
		12'd 2567 : data_o = 23'b 10000010111110001111110 ;
		12'd 2568 : data_o = 23'b 10000010110110110100001 ;
		12'd 2569 : data_o = 23'b 10000010101111011000101 ;
		12'd 2570 : data_o = 23'b 10000010100111111101011 ;
		12'd 2571 : data_o = 23'b 10000010100000100010011 ;
		12'd 2572 : data_o = 23'b 10000010011001000111100 ;
		12'd 2573 : data_o = 23'b 10000010010001101101000 ;
		12'd 2574 : data_o = 23'b 10000010001010010010101 ;
		12'd 2575 : data_o = 23'b 10000010000010111000011 ;
		12'd 2576 : data_o = 23'b 10000001111011011110100 ;
		12'd 2577 : data_o = 23'b 10000001110100000100110 ;
		12'd 2578 : data_o = 23'b 10000001101100101011001 ;
		12'd 2579 : data_o = 23'b 10000001100101010001111 ;
		12'd 2580 : data_o = 23'b 10000001011101111000110 ;
		12'd 2581 : data_o = 23'b 10000001010110011111111 ;
		12'd 2582 : data_o = 23'b 10000001001111000111001 ;
		12'd 2583 : data_o = 23'b 10000001000111101110110 ;
		12'd 2584 : data_o = 23'b 10000001000000010110100 ;
		12'd 2585 : data_o = 23'b 10000000111000111110011 ;
		12'd 2586 : data_o = 23'b 10000000110001100110101 ;
		12'd 2587 : data_o = 23'b 10000000101010001111000 ;
		12'd 2588 : data_o = 23'b 10000000100010110111100 ;
		12'd 2589 : data_o = 23'b 10000000011011100000011 ;
		12'd 2590 : data_o = 23'b 10000000010100001001011 ;
		12'd 2591 : data_o = 23'b 10000000001100110010101 ;
		12'd 2592 : data_o = 23'b 10000000000101011100000 ;
		12'd 2593 : data_o = 23'b 01111111111110000101101 ;
		12'd 2594 : data_o = 23'b 01111111110110101111100 ;
		12'd 2595 : data_o = 23'b 01111111101111011001101 ;
		12'd 2596 : data_o = 23'b 01111111101000000011111 ;
		12'd 2597 : data_o = 23'b 01111111100000101110011 ;
		12'd 2598 : data_o = 23'b 01111111011001011001000 ;
		12'd 2599 : data_o = 23'b 01111111010010000100000 ;
		12'd 2600 : data_o = 23'b 01111111001010101111001 ;
		12'd 2601 : data_o = 23'b 01111111000011011010011 ;
		12'd 2602 : data_o = 23'b 01111110111100000110000 ;
		12'd 2603 : data_o = 23'b 01111110110100110001110 ;
		12'd 2604 : data_o = 23'b 01111110101101011101101 ;
		12'd 2605 : data_o = 23'b 01111110100110001001111 ;
		12'd 2606 : data_o = 23'b 01111110011110110110010 ;
		12'd 2607 : data_o = 23'b 01111110010111100010111 ;
		12'd 2608 : data_o = 23'b 01111110010000001111101 ;
		12'd 2609 : data_o = 23'b 01111110001000111100101 ;
		12'd 2610 : data_o = 23'b 01111110000001101001111 ;
		12'd 2611 : data_o = 23'b 01111101111010010111010 ;
		12'd 2612 : data_o = 23'b 01111101110011000100111 ;
		12'd 2613 : data_o = 23'b 01111101101011110010110 ;
		12'd 2614 : data_o = 23'b 01111101100100100000110 ;
		12'd 2615 : data_o = 23'b 01111101011101001111000 ;
		12'd 2616 : data_o = 23'b 01111101010101111101100 ;
		12'd 2617 : data_o = 23'b 01111101001110101100001 ;
		12'd 2618 : data_o = 23'b 01111101000111011011001 ;
		12'd 2619 : data_o = 23'b 01111101000000001010001 ;
		12'd 2620 : data_o = 23'b 01111100111000111001100 ;
		12'd 2621 : data_o = 23'b 01111100110001101001000 ;
		12'd 2622 : data_o = 23'b 01111100101010011000101 ;
		12'd 2623 : data_o = 23'b 01111100100011001000101 ;
		12'd 2624 : data_o = 23'b 01111100011011111000110 ;
		12'd 2625 : data_o = 23'b 01111100010100101001000 ;
		12'd 2626 : data_o = 23'b 01111100001101011001101 ;
		12'd 2627 : data_o = 23'b 01111100000110001010011 ;
		12'd 2628 : data_o = 23'b 01111011111110111011010 ;
		12'd 2629 : data_o = 23'b 01111011110111101100100 ;
		12'd 2630 : data_o = 23'b 01111011110000011101111 ;
		12'd 2631 : data_o = 23'b 01111011101001001111011 ;
		12'd 2632 : data_o = 23'b 01111011100010000001001 ;
		12'd 2633 : data_o = 23'b 01111011011010110011001 ;
		12'd 2634 : data_o = 23'b 01111011010011100101011 ;
		12'd 2635 : data_o = 23'b 01111011001100010111110 ;
		12'd 2636 : data_o = 23'b 01111011000101001010011 ;
		12'd 2637 : data_o = 23'b 01111010111101111101001 ;
		12'd 2638 : data_o = 23'b 01111010110110110000001 ;
		12'd 2639 : data_o = 23'b 01111010101111100011011 ;
		12'd 2640 : data_o = 23'b 01111010101000010110111 ;
		12'd 2641 : data_o = 23'b 01111010100001001010100 ;
		12'd 2642 : data_o = 23'b 01111010011001111110010 ;
		12'd 2643 : data_o = 23'b 01111010010010110010011 ;
		12'd 2644 : data_o = 23'b 01111010001011100110101 ;
		12'd 2645 : data_o = 23'b 01111010000100011011000 ;
		12'd 2646 : data_o = 23'b 01111001111101001111101 ;
		12'd 2647 : data_o = 23'b 01111001110110000100100 ;
		12'd 2648 : data_o = 23'b 01111001101110111001101 ;
		12'd 2649 : data_o = 23'b 01111001100111101110111 ;
		12'd 2650 : data_o = 23'b 01111001100000100100011 ;
		12'd 2651 : data_o = 23'b 01111001011001011010000 ;
		12'd 2652 : data_o = 23'b 01111001010010001111111 ;
		12'd 2653 : data_o = 23'b 01111001001011000110000 ;
		12'd 2654 : data_o = 23'b 01111001000011111100010 ;
		12'd 2655 : data_o = 23'b 01111000111100110010110 ;
		12'd 2656 : data_o = 23'b 01111000110101101001011 ;
		12'd 2657 : data_o = 23'b 01111000101110100000011 ;
		12'd 2658 : data_o = 23'b 01111000100111010111011 ;
		12'd 2659 : data_o = 23'b 01111000100000001110110 ;
		12'd 2660 : data_o = 23'b 01111000011001000110010 ;
		12'd 2661 : data_o = 23'b 01111000010001111110000 ;
		12'd 2662 : data_o = 23'b 01111000001010110101111 ;
		12'd 2663 : data_o = 23'b 01111000000011101110000 ;
		12'd 2664 : data_o = 23'b 01110111111100100110010 ;
		12'd 2665 : data_o = 23'b 01110111110101011110110 ;
		12'd 2666 : data_o = 23'b 01110111101110010111100 ;
		12'd 2667 : data_o = 23'b 01110111100111010000011 ;
		12'd 2668 : data_o = 23'b 01110111100000001001100 ;
		12'd 2669 : data_o = 23'b 01110111011001000010111 ;
		12'd 2670 : data_o = 23'b 01110111010001111100011 ;
		12'd 2671 : data_o = 23'b 01110111001010110110001 ;
		12'd 2672 : data_o = 23'b 01110111000011110000000 ;
		12'd 2673 : data_o = 23'b 01110110111100101010001 ;
		12'd 2674 : data_o = 23'b 01110110110101100100100 ;
		12'd 2675 : data_o = 23'b 01110110101110011111000 ;
		12'd 2676 : data_o = 23'b 01110110100111011001110 ;
		12'd 2677 : data_o = 23'b 01110110100000010100110 ;
		12'd 2678 : data_o = 23'b 01110110011001001111111 ;
		12'd 2679 : data_o = 23'b 01110110010010001011001 ;
		12'd 2680 : data_o = 23'b 01110110001011000110110 ;
		12'd 2681 : data_o = 23'b 01110110000100000010100 ;
		12'd 2682 : data_o = 23'b 01110101111100111110011 ;
		12'd 2683 : data_o = 23'b 01110101110101111010100 ;
		12'd 2684 : data_o = 23'b 01110101101110110110111 ;
		12'd 2685 : data_o = 23'b 01110101100111110011011 ;
		12'd 2686 : data_o = 23'b 01110101100000110000001 ;
		12'd 2687 : data_o = 23'b 01110101011001101101000 ;
		12'd 2688 : data_o = 23'b 01110101010010101010001 ;
		12'd 2689 : data_o = 23'b 01110101001011100111100 ;
		12'd 2690 : data_o = 23'b 01110101000100100101000 ;
		12'd 2691 : data_o = 23'b 01110100111101100010110 ;
		12'd 2692 : data_o = 23'b 01110100110110100000110 ;
		12'd 2693 : data_o = 23'b 01110100101111011110111 ;
		12'd 2694 : data_o = 23'b 01110100101000011101001 ;
		12'd 2695 : data_o = 23'b 01110100100001011011101 ;
		12'd 2696 : data_o = 23'b 01110100011010011010011 ;
		12'd 2697 : data_o = 23'b 01110100010011011001011 ;
		12'd 2698 : data_o = 23'b 01110100001100011000100 ;
		12'd 2699 : data_o = 23'b 01110100000101010111110 ;
		12'd 2700 : data_o = 23'b 01110011111110010111010 ;
		12'd 2701 : data_o = 23'b 01110011110111010111000 ;
		12'd 2702 : data_o = 23'b 01110011110000010110111 ;
		12'd 2703 : data_o = 23'b 01110011101001010111000 ;
		12'd 2704 : data_o = 23'b 01110011100010010111011 ;
		12'd 2705 : data_o = 23'b 01110011011011010111111 ;
		12'd 2706 : data_o = 23'b 01110011010100011000100 ;
		12'd 2707 : data_o = 23'b 01110011001101011001100 ;
		12'd 2708 : data_o = 23'b 01110011000110011010100 ;
		12'd 2709 : data_o = 23'b 01110010111111011011111 ;
		12'd 2710 : data_o = 23'b 01110010111000011101011 ;
		12'd 2711 : data_o = 23'b 01110010110001011111000 ;
		12'd 2712 : data_o = 23'b 01110010101010100000111 ;
		12'd 2713 : data_o = 23'b 01110010100011100011000 ;
		12'd 2714 : data_o = 23'b 01110010011100100101010 ;
		12'd 2715 : data_o = 23'b 01110010010101100111110 ;
		12'd 2716 : data_o = 23'b 01110010001110101010011 ;
		12'd 2717 : data_o = 23'b 01110010000111101101010 ;
		12'd 2718 : data_o = 23'b 01110010000000110000011 ;
		12'd 2719 : data_o = 23'b 01110001111001110011101 ;
		12'd 2720 : data_o = 23'b 01110001110010110111000 ;
		12'd 2721 : data_o = 23'b 01110001101011111010110 ;
		12'd 2722 : data_o = 23'b 01110001100100111110100 ;
		12'd 2723 : data_o = 23'b 01110001011110000010101 ;
		12'd 2724 : data_o = 23'b 01110001010111000110111 ;
		12'd 2725 : data_o = 23'b 01110001010000001011010 ;
		12'd 2726 : data_o = 23'b 01110001001001001111111 ;
		12'd 2727 : data_o = 23'b 01110001000010010100110 ;
		12'd 2728 : data_o = 23'b 01110000111011011001110 ;
		12'd 2729 : data_o = 23'b 01110000110100011110111 ;
		12'd 2730 : data_o = 23'b 01110000101101100100011 ;
		12'd 2731 : data_o = 23'b 01110000100110101001111 ;
		12'd 2732 : data_o = 23'b 01110000011111101111110 ;
		12'd 2733 : data_o = 23'b 01110000011000110101110 ;
		12'd 2734 : data_o = 23'b 01110000010001111011111 ;
		12'd 2735 : data_o = 23'b 01110000001011000010010 ;
		12'd 2736 : data_o = 23'b 01110000000100001000111 ;
		12'd 2737 : data_o = 23'b 01101111111101001111101 ;
		12'd 2738 : data_o = 23'b 01101111110110010110101 ;
		12'd 2739 : data_o = 23'b 01101111101111011101110 ;
		12'd 2740 : data_o = 23'b 01101111101000100101000 ;
		12'd 2741 : data_o = 23'b 01101111100001101100101 ;
		12'd 2742 : data_o = 23'b 01101111011010110100011 ;
		12'd 2743 : data_o = 23'b 01101111010011111100010 ;
		12'd 2744 : data_o = 23'b 01101111001101000100011 ;
		12'd 2745 : data_o = 23'b 01101111000110001100101 ;
		12'd 2746 : data_o = 23'b 01101110111111010101001 ;
		12'd 2747 : data_o = 23'b 01101110111000011101111 ;
		12'd 2748 : data_o = 23'b 01101110110001100110110 ;
		12'd 2749 : data_o = 23'b 01101110101010101111111 ;
		12'd 2750 : data_o = 23'b 01101110100011111001001 ;
		12'd 2751 : data_o = 23'b 01101110011101000010101 ;
		12'd 2752 : data_o = 23'b 01101110010110001100010 ;
		12'd 2753 : data_o = 23'b 01101110001111010110001 ;
		12'd 2754 : data_o = 23'b 01101110001000100000001 ;
		12'd 2755 : data_o = 23'b 01101110000001101010011 ;
		12'd 2756 : data_o = 23'b 01101101111010110100110 ;
		12'd 2757 : data_o = 23'b 01101101110011111111011 ;
		12'd 2758 : data_o = 23'b 01101101101101001010010 ;
		12'd 2759 : data_o = 23'b 01101101100110010101010 ;
		12'd 2760 : data_o = 23'b 01101101011111100000011 ;
		12'd 2761 : data_o = 23'b 01101101011000101011110 ;
		12'd 2762 : data_o = 23'b 01101101010001110111011 ;
		12'd 2763 : data_o = 23'b 01101101001011000011001 ;
		12'd 2764 : data_o = 23'b 01101101000100001111001 ;
		12'd 2765 : data_o = 23'b 01101100111101011011010 ;
		12'd 2766 : data_o = 23'b 01101100110110100111100 ;
		12'd 2767 : data_o = 23'b 01101100101111110100001 ;
		12'd 2768 : data_o = 23'b 01101100101001000000110 ;
		12'd 2769 : data_o = 23'b 01101100100010001101110 ;
		12'd 2770 : data_o = 23'b 01101100011011011010110 ;
		12'd 2771 : data_o = 23'b 01101100010100101000001 ;
		12'd 2772 : data_o = 23'b 01101100001101110101101 ;
		12'd 2773 : data_o = 23'b 01101100000111000011010 ;
		12'd 2774 : data_o = 23'b 01101100000000010001001 ;
		12'd 2775 : data_o = 23'b 01101011111001011111001 ;
		12'd 2776 : data_o = 23'b 01101011110010101101011 ;
		12'd 2777 : data_o = 23'b 01101011101011111011110 ;
		12'd 2778 : data_o = 23'b 01101011100101001010011 ;
		12'd 2779 : data_o = 23'b 01101011011110011001010 ;
		12'd 2780 : data_o = 23'b 01101011010111101000010 ;
		12'd 2781 : data_o = 23'b 01101011010000110111011 ;
		12'd 2782 : data_o = 23'b 01101011001010000110110 ;
		12'd 2783 : data_o = 23'b 01101011000011010110010 ;
		12'd 2784 : data_o = 23'b 01101010111100100110000 ;
		12'd 2785 : data_o = 23'b 01101010110101110110000 ;
		12'd 2786 : data_o = 23'b 01101010101111000110001 ;
		12'd 2787 : data_o = 23'b 01101010101000010110011 ;
		12'd 2788 : data_o = 23'b 01101010100001100110111 ;
		12'd 2789 : data_o = 23'b 01101010011010110111101 ;
		12'd 2790 : data_o = 23'b 01101010010100001000100 ;
		12'd 2791 : data_o = 23'b 01101010001101011001100 ;
		12'd 2792 : data_o = 23'b 01101010000110101010110 ;
		12'd 2793 : data_o = 23'b 01101001111111111100010 ;
		12'd 2794 : data_o = 23'b 01101001111001001101111 ;
		12'd 2795 : data_o = 23'b 01101001110010011111101 ;
		12'd 2796 : data_o = 23'b 01101001101011110001101 ;
		12'd 2797 : data_o = 23'b 01101001100101000011111 ;
		12'd 2798 : data_o = 23'b 01101001011110010110010 ;
		12'd 2799 : data_o = 23'b 01101001010111101000110 ;
		12'd 2800 : data_o = 23'b 01101001010000111011100 ;
		12'd 2801 : data_o = 23'b 01101001001010001110100 ;
		12'd 2802 : data_o = 23'b 01101001000011100001101 ;
		12'd 2803 : data_o = 23'b 01101000111100110100111 ;
		12'd 2804 : data_o = 23'b 01101000110110001000011 ;
		12'd 2805 : data_o = 23'b 01101000101111011100001 ;
		12'd 2806 : data_o = 23'b 01101000101000101111111 ;
		12'd 2807 : data_o = 23'b 01101000100010000100000 ;
		12'd 2808 : data_o = 23'b 01101000011011011000010 ;
		12'd 2809 : data_o = 23'b 01101000010100101100101 ;
		12'd 2810 : data_o = 23'b 01101000001110000001010 ;
		12'd 2811 : data_o = 23'b 01101000000111010110000 ;
		12'd 2812 : data_o = 23'b 01101000000000101011000 ;
		12'd 2813 : data_o = 23'b 01100111111010000000010 ;
		12'd 2814 : data_o = 23'b 01100111110011010101100 ;
		12'd 2815 : data_o = 23'b 01100111101100101011001 ;
		12'd 2816 : data_o = 23'b 01100111100110000000111 ;
		12'd 2817 : data_o = 23'b 01100111011111010110110 ;
		12'd 2818 : data_o = 23'b 01100111011000101100111 ;
		12'd 2819 : data_o = 23'b 01100111010010000011001 ;
		12'd 2820 : data_o = 23'b 01100111001011011001100 ;
		12'd 2821 : data_o = 23'b 01100111000100110000010 ;
		12'd 2822 : data_o = 23'b 01100110111110000111000 ;
		12'd 2823 : data_o = 23'b 01100110110111011110000 ;
		12'd 2824 : data_o = 23'b 01100110110000110101010 ;
		12'd 2825 : data_o = 23'b 01100110101010001100101 ;
		12'd 2826 : data_o = 23'b 01100110100011100100010 ;
		12'd 2827 : data_o = 23'b 01100110011100111100000 ;
		12'd 2828 : data_o = 23'b 01100110010110010011111 ;
		12'd 2829 : data_o = 23'b 01100110001111101100000 ;
		12'd 2830 : data_o = 23'b 01100110001001000100010 ;
		12'd 2831 : data_o = 23'b 01100110000010011100110 ;
		12'd 2832 : data_o = 23'b 01100101111011110101100 ;
		12'd 2833 : data_o = 23'b 01100101110101001110010 ;
		12'd 2834 : data_o = 23'b 01100101101110100111011 ;
		12'd 2835 : data_o = 23'b 01100101101000000000100 ;
		12'd 2836 : data_o = 23'b 01100101100001011010000 ;
		12'd 2837 : data_o = 23'b 01100101011010110011100 ;
		12'd 2838 : data_o = 23'b 01100101010100001101010 ;
		12'd 2839 : data_o = 23'b 01100101001101100111010 ;
		12'd 2840 : data_o = 23'b 01100101000111000001011 ;
		12'd 2841 : data_o = 23'b 01100101000000011011110 ;
		12'd 2842 : data_o = 23'b 01100100111001110110010 ;
		12'd 2843 : data_o = 23'b 01100100110011010000111 ;
		12'd 2844 : data_o = 23'b 01100100101100101011110 ;
		12'd 2845 : data_o = 23'b 01100100100110000110110 ;
		12'd 2846 : data_o = 23'b 01100100011111100010000 ;
		12'd 2847 : data_o = 23'b 01100100011000111101011 ;
		12'd 2848 : data_o = 23'b 01100100010010011001000 ;
		12'd 2849 : data_o = 23'b 01100100001011110100110 ;
		12'd 2850 : data_o = 23'b 01100100000101010000110 ;
		12'd 2851 : data_o = 23'b 01100011111110101100111 ;
		12'd 2852 : data_o = 23'b 01100011111000001001001 ;
		12'd 2853 : data_o = 23'b 01100011110001100101101 ;
		12'd 2854 : data_o = 23'b 01100011101011000010011 ;
		12'd 2855 : data_o = 23'b 01100011100100011111010 ;
		12'd 2856 : data_o = 23'b 01100011011101111100010 ;
		12'd 2857 : data_o = 23'b 01100011010111011001100 ;
		12'd 2858 : data_o = 23'b 01100011010000110110111 ;
		12'd 2859 : data_o = 23'b 01100011001010010100100 ;
		12'd 2860 : data_o = 23'b 01100011000011110010010 ;
		12'd 2861 : data_o = 23'b 01100010111101010000001 ;
		12'd 2862 : data_o = 23'b 01100010110110101110010 ;
		12'd 2863 : data_o = 23'b 01100010110000001100101 ;
		12'd 2864 : data_o = 23'b 01100010101001101011000 ;
		12'd 2865 : data_o = 23'b 01100010100011001001110 ;
		12'd 2866 : data_o = 23'b 01100010011100101000100 ;
		12'd 2867 : data_o = 23'b 01100010010110000111101 ;
		12'd 2868 : data_o = 23'b 01100010001111100110110 ;
		12'd 2869 : data_o = 23'b 01100010001001000110001 ;
		12'd 2870 : data_o = 23'b 01100010000010100101110 ;
		12'd 2871 : data_o = 23'b 01100001111100000101100 ;
		12'd 2872 : data_o = 23'b 01100001110101100101011 ;
		12'd 2873 : data_o = 23'b 01100001101111000101100 ;
		12'd 2874 : data_o = 23'b 01100001101000100101110 ;
		12'd 2875 : data_o = 23'b 01100001100010000110010 ;
		12'd 2876 : data_o = 23'b 01100001011011100110111 ;
		12'd 2877 : data_o = 23'b 01100001010101000111101 ;
		12'd 2878 : data_o = 23'b 01100001001110101000101 ;
		12'd 2879 : data_o = 23'b 01100001001000001001110 ;
		12'd 2880 : data_o = 23'b 01100001000001101011001 ;
		12'd 2881 : data_o = 23'b 01100000111011001100101 ;
		12'd 2882 : data_o = 23'b 01100000110100101110011 ;
		12'd 2883 : data_o = 23'b 01100000101110010000010 ;
		12'd 2884 : data_o = 23'b 01100000100111110010011 ;
		12'd 2885 : data_o = 23'b 01100000100001010100101 ;
		12'd 2886 : data_o = 23'b 01100000011010110111000 ;
		12'd 2887 : data_o = 23'b 01100000010100011001101 ;
		12'd 2888 : data_o = 23'b 01100000001101111100011 ;
		12'd 2889 : data_o = 23'b 01100000000111011111010 ;
		12'd 2890 : data_o = 23'b 01100000000001000010011 ;
		12'd 2891 : data_o = 23'b 01011111111010100101110 ;
		12'd 2892 : data_o = 23'b 01011111110100001001010 ;
		12'd 2893 : data_o = 23'b 01011111101101101100111 ;
		12'd 2894 : data_o = 23'b 01011111100111010000110 ;
		12'd 2895 : data_o = 23'b 01011111100000110100110 ;
		12'd 2896 : data_o = 23'b 01011111011010011000111 ;
		12'd 2897 : data_o = 23'b 01011111010011111101010 ;
		12'd 2898 : data_o = 23'b 01011111001101100001110 ;
		12'd 2899 : data_o = 23'b 01011111000111000110100 ;
		12'd 2900 : data_o = 23'b 01011111000000101011011 ;
		12'd 2901 : data_o = 23'b 01011110111010010000100 ;
		12'd 2902 : data_o = 23'b 01011110110011110101110 ;
		12'd 2903 : data_o = 23'b 01011110101101011011001 ;
		12'd 2904 : data_o = 23'b 01011110100111000000110 ;
		12'd 2905 : data_o = 23'b 01011110100000100110100 ;
		12'd 2906 : data_o = 23'b 01011110011010001100100 ;
		12'd 2907 : data_o = 23'b 01011110010011110010101 ;
		12'd 2908 : data_o = 23'b 01011110001101011000111 ;
		12'd 2909 : data_o = 23'b 01011110000110111111011 ;
		12'd 2910 : data_o = 23'b 01011110000000100110000 ;
		12'd 2911 : data_o = 23'b 01011101111010001100111 ;
		12'd 2912 : data_o = 23'b 01011101110011110011111 ;
		12'd 2913 : data_o = 23'b 01011101101101011011000 ;
		12'd 2914 : data_o = 23'b 01011101100111000010011 ;
		12'd 2915 : data_o = 23'b 01011101100000101001111 ;
		12'd 2916 : data_o = 23'b 01011101011010010001101 ;
		12'd 2917 : data_o = 23'b 01011101010011111001100 ;
		12'd 2918 : data_o = 23'b 01011101001101100001100 ;
		12'd 2919 : data_o = 23'b 01011101000111001001110 ;
		12'd 2920 : data_o = 23'b 01011101000000110010001 ;
		12'd 2921 : data_o = 23'b 01011100111010011010110 ;
		12'd 2922 : data_o = 23'b 01011100110100000011100 ;
		12'd 2923 : data_o = 23'b 01011100101101101100011 ;
		12'd 2924 : data_o = 23'b 01011100100111010101100 ;
		12'd 2925 : data_o = 23'b 01011100100000111110110 ;
		12'd 2926 : data_o = 23'b 01011100011010101000010 ;
		12'd 2927 : data_o = 23'b 01011100010100010001111 ;
		12'd 2928 : data_o = 23'b 01011100001101111011101 ;
		12'd 2929 : data_o = 23'b 01011100000111100101101 ;
		12'd 2930 : data_o = 23'b 01011100000001001111110 ;
		12'd 2931 : data_o = 23'b 01011011111010111010001 ;
		12'd 2932 : data_o = 23'b 01011011110100100100100 ;
		12'd 2933 : data_o = 23'b 01011011101110001111010 ;
		12'd 2934 : data_o = 23'b 01011011100111111010000 ;
		12'd 2935 : data_o = 23'b 01011011100001100101000 ;
		12'd 2936 : data_o = 23'b 01011011011011010000010 ;
		12'd 2937 : data_o = 23'b 01011011010100111011101 ;
		12'd 2938 : data_o = 23'b 01011011001110100111001 ;
		12'd 2939 : data_o = 23'b 01011011001000010010110 ;
		12'd 2940 : data_o = 23'b 01011011000001111110101 ;
		12'd 2941 : data_o = 23'b 01011010111011101010110 ;
		12'd 2942 : data_o = 23'b 01011010110101010110111 ;
		12'd 2943 : data_o = 23'b 01011010101111000011010 ;
		12'd 2944 : data_o = 23'b 01011010101000101111111 ;
		12'd 2945 : data_o = 23'b 01011010100010011100101 ;
		12'd 2946 : data_o = 23'b 01011010011100001001100 ;
		12'd 2947 : data_o = 23'b 01011010010101110110100 ;
		12'd 2948 : data_o = 23'b 01011010001111100011110 ;
		12'd 2949 : data_o = 23'b 01011010001001010001010 ;
		12'd 2950 : data_o = 23'b 01011010000010111110110 ;
		12'd 2951 : data_o = 23'b 01011001111100101100100 ;
		12'd 2952 : data_o = 23'b 01011001110110011010100 ;
		12'd 2953 : data_o = 23'b 01011001110000001000100 ;
		12'd 2954 : data_o = 23'b 01011001101001110110111 ;
		12'd 2955 : data_o = 23'b 01011001100011100101010 ;
		12'd 2956 : data_o = 23'b 01011001011101010011111 ;
		12'd 2957 : data_o = 23'b 01011001010111000010101 ;
		12'd 2958 : data_o = 23'b 01011001010000110001101 ;
		12'd 2959 : data_o = 23'b 01011001001010100000110 ;
		12'd 2960 : data_o = 23'b 01011001000100010000000 ;
		12'd 2961 : data_o = 23'b 01011000111101111111100 ;
		12'd 2962 : data_o = 23'b 01011000110111101111001 ;
		12'd 2963 : data_o = 23'b 01011000110001011110111 ;
		12'd 2964 : data_o = 23'b 01011000101011001110111 ;
		12'd 2965 : data_o = 23'b 01011000100100111111000 ;
		12'd 2966 : data_o = 23'b 01011000011110101111011 ;
		12'd 2967 : data_o = 23'b 01011000011000011111111 ;
		12'd 2968 : data_o = 23'b 01011000010010010000100 ;
		12'd 2969 : data_o = 23'b 01011000001100000001011 ;
		12'd 2970 : data_o = 23'b 01011000000101110010011 ;
		12'd 2971 : data_o = 23'b 01010111111111100011100 ;
		12'd 2972 : data_o = 23'b 01010111111001010100110 ;
		12'd 2973 : data_o = 23'b 01010111110011000110010 ;
		12'd 2974 : data_o = 23'b 01010111101100111000000 ;
		12'd 2975 : data_o = 23'b 01010111100110101001111 ;
		12'd 2976 : data_o = 23'b 01010111100000011011111 ;
		12'd 2977 : data_o = 23'b 01010111011010001110000 ;
		12'd 2978 : data_o = 23'b 01010111010100000000011 ;
		12'd 2979 : data_o = 23'b 01010111001101110010111 ;
		12'd 2980 : data_o = 23'b 01010111000111100101100 ;
		12'd 2981 : data_o = 23'b 01010111000001011000011 ;
		12'd 2982 : data_o = 23'b 01010110111011001011011 ;
		12'd 2983 : data_o = 23'b 01010110110100111110101 ;
		12'd 2984 : data_o = 23'b 01010110101110110010000 ;
		12'd 2985 : data_o = 23'b 01010110101000100101100 ;
		12'd 2986 : data_o = 23'b 01010110100010011001001 ;
		12'd 2987 : data_o = 23'b 01010110011100001101000 ;
		12'd 2988 : data_o = 23'b 01010110010110000001000 ;
		12'd 2989 : data_o = 23'b 01010110001111110101010 ;
		12'd 2990 : data_o = 23'b 01010110001001101001101 ;
		12'd 2991 : data_o = 23'b 01010110000011011110001 ;
		12'd 2992 : data_o = 23'b 01010101111101010010111 ;
		12'd 2993 : data_o = 23'b 01010101110111000111110 ;
		12'd 2994 : data_o = 23'b 01010101110000111100110 ;
		12'd 2995 : data_o = 23'b 01010101101010110001111 ;
		12'd 2996 : data_o = 23'b 01010101100100100111010 ;
		12'd 2997 : data_o = 23'b 01010101011110011100111 ;
		12'd 2998 : data_o = 23'b 01010101011000010010100 ;
		12'd 2999 : data_o = 23'b 01010101010010001000011 ;
		12'd 3000 : data_o = 23'b 01010101001011111110011 ;
		12'd 3001 : data_o = 23'b 01010101000101110100101 ;
		12'd 3002 : data_o = 23'b 01010100111111101011000 ;
		12'd 3003 : data_o = 23'b 01010100111001100001100 ;
		12'd 3004 : data_o = 23'b 01010100110011011000010 ;
		12'd 3005 : data_o = 23'b 01010100101101001111001 ;
		12'd 3006 : data_o = 23'b 01010100100111000110001 ;
		12'd 3007 : data_o = 23'b 01010100100000111101010 ;
		12'd 3008 : data_o = 23'b 01010100011010110100101 ;
		12'd 3009 : data_o = 23'b 01010100010100101100010 ;
		12'd 3010 : data_o = 23'b 01010100001110100011111 ;
		12'd 3011 : data_o = 23'b 01010100001000011011110 ;
		12'd 3012 : data_o = 23'b 01010100000010010011110 ;
		12'd 3013 : data_o = 23'b 01010011111100001100000 ;
		12'd 3014 : data_o = 23'b 01010011110110000100010 ;
		12'd 3015 : data_o = 23'b 01010011101111111100111 ;
		12'd 3016 : data_o = 23'b 01010011101001110101100 ;
		12'd 3017 : data_o = 23'b 01010011100011101110011 ;
		12'd 3018 : data_o = 23'b 01010011011101100111011 ;
		12'd 3019 : data_o = 23'b 01010011010111100000100 ;
		12'd 3020 : data_o = 23'b 01010011010001011001111 ;
		12'd 3021 : data_o = 23'b 01010011001011010011011 ;
		12'd 3022 : data_o = 23'b 01010011000101001101001 ;
		12'd 3023 : data_o = 23'b 01010010111111000110111 ;
		12'd 3024 : data_o = 23'b 01010010111001000000111 ;
		12'd 3025 : data_o = 23'b 01010010110010111011001 ;
		12'd 3026 : data_o = 23'b 01010010101100110101011 ;
		12'd 3027 : data_o = 23'b 01010010100110101111111 ;
		12'd 3028 : data_o = 23'b 01010010100000101010101 ;
		12'd 3029 : data_o = 23'b 01010010011010100101011 ;
		12'd 3030 : data_o = 23'b 01010010010100100000011 ;
		12'd 3031 : data_o = 23'b 01010010001110011011100 ;
		12'd 3032 : data_o = 23'b 01010010001000010110111 ;
		12'd 3033 : data_o = 23'b 01010010000010010010011 ;
		12'd 3034 : data_o = 23'b 01010001111100001110000 ;
		12'd 3035 : data_o = 23'b 01010001110110001001110 ;
		12'd 3036 : data_o = 23'b 01010001110000000101110 ;
		12'd 3037 : data_o = 23'b 01010001101010000001111 ;
		12'd 3038 : data_o = 23'b 01010001100011111110001 ;
		12'd 3039 : data_o = 23'b 01010001011101111010101 ;
		12'd 3040 : data_o = 23'b 01010001010111110111010 ;
		12'd 3041 : data_o = 23'b 01010001010001110100000 ;
		12'd 3042 : data_o = 23'b 01010001001011110001000 ;
		12'd 3043 : data_o = 23'b 01010001000101101110001 ;
		12'd 3044 : data_o = 23'b 01010000111111101011011 ;
		12'd 3045 : data_o = 23'b 01010000111001101000110 ;
		12'd 3046 : data_o = 23'b 01010000110011100110011 ;
		12'd 3047 : data_o = 23'b 01010000101101100100001 ;
		12'd 3048 : data_o = 23'b 01010000100111100010001 ;
		12'd 3049 : data_o = 23'b 01010000100001100000001 ;
		12'd 3050 : data_o = 23'b 01010000011011011110011 ;
		12'd 3051 : data_o = 23'b 01010000010101011100110 ;
		12'd 3052 : data_o = 23'b 01010000001111011011011 ;
		12'd 3053 : data_o = 23'b 01010000001001011010001 ;
		12'd 3054 : data_o = 23'b 01010000000011011001000 ;
		12'd 3055 : data_o = 23'b 01001111111101011000000 ;
		12'd 3056 : data_o = 23'b 01001111110111010111010 ;
		12'd 3057 : data_o = 23'b 01001111110001010110101 ;
		12'd 3058 : data_o = 23'b 01001111101011010110001 ;
		12'd 3059 : data_o = 23'b 01001111100101010101111 ;
		12'd 3060 : data_o = 23'b 01001111011111010101110 ;
		12'd 3061 : data_o = 23'b 01001111011001010101110 ;
		12'd 3062 : data_o = 23'b 01001111010011010110000 ;
		12'd 3063 : data_o = 23'b 01001111001101010110010 ;
		12'd 3064 : data_o = 23'b 01001111000111010110110 ;
		12'd 3065 : data_o = 23'b 01001111000001010111100 ;
		12'd 3066 : data_o = 23'b 01001110111011011000010 ;
		12'd 3067 : data_o = 23'b 01001110110101011001010 ;
		12'd 3068 : data_o = 23'b 01001110101111011010011 ;
		12'd 3069 : data_o = 23'b 01001110101001011011110 ;
		12'd 3070 : data_o = 23'b 01001110100011011101001 ;
		12'd 3071 : data_o = 23'b 01001110011101011110110 ;
		12'd 3072 : data_o = 23'b 01001110010111100000101 ;
		12'd 3073 : data_o = 23'b 01001110010001100010100 ;
		12'd 3074 : data_o = 23'b 01001110001011100100101 ;
		12'd 3075 : data_o = 23'b 01001110000101100110111 ;
		12'd 3076 : data_o = 23'b 01001101111111101001011 ;
		12'd 3077 : data_o = 23'b 01001101111001101011111 ;
		12'd 3078 : data_o = 23'b 01001101110011101110101 ;
		12'd 3079 : data_o = 23'b 01001101101101110001101 ;
		12'd 3080 : data_o = 23'b 01001101100111110100101 ;
		12'd 3081 : data_o = 23'b 01001101100001110111111 ;
		12'd 3082 : data_o = 23'b 01001101011011111011010 ;
		12'd 3083 : data_o = 23'b 01001101010101111110110 ;
		12'd 3084 : data_o = 23'b 01001101010000000010100 ;
		12'd 3085 : data_o = 23'b 01001101001010000110011 ;
		12'd 3086 : data_o = 23'b 01001101000100001010011 ;
		12'd 3087 : data_o = 23'b 01001100111110001110100 ;
		12'd 3088 : data_o = 23'b 01001100111000010010111 ;
		12'd 3089 : data_o = 23'b 01001100110010010111011 ;
		12'd 3090 : data_o = 23'b 01001100101100011100000 ;
		12'd 3091 : data_o = 23'b 01001100100110100000110 ;
		12'd 3092 : data_o = 23'b 01001100100000100101110 ;
		12'd 3093 : data_o = 23'b 01001100011010101010111 ;
		12'd 3094 : data_o = 23'b 01001100010100110000001 ;
		12'd 3095 : data_o = 23'b 01001100001110110101101 ;
		12'd 3096 : data_o = 23'b 01001100001000111011010 ;
		12'd 3097 : data_o = 23'b 01001100000011000001000 ;
		12'd 3098 : data_o = 23'b 01001011111101000110111 ;
		12'd 3099 : data_o = 23'b 01001011110111001101000 ;
		12'd 3100 : data_o = 23'b 01001011110001010011010 ;
		12'd 3101 : data_o = 23'b 01001011101011011001101 ;
		12'd 3102 : data_o = 23'b 01001011100101100000001 ;
		12'd 3103 : data_o = 23'b 01001011011111100110111 ;
		12'd 3104 : data_o = 23'b 01001011011001101101110 ;
		12'd 3105 : data_o = 23'b 01001011010011110100110 ;
		12'd 3106 : data_o = 23'b 01001011001101111011111 ;
		12'd 3107 : data_o = 23'b 01001011001000000011010 ;
		12'd 3108 : data_o = 23'b 01001011000010001010110 ;
		12'd 3109 : data_o = 23'b 01001010111100010010011 ;
		12'd 3110 : data_o = 23'b 01001010110110011010001 ;
		12'd 3111 : data_o = 23'b 01001010110000100010001 ;
		12'd 3112 : data_o = 23'b 01001010101010101010010 ;
		12'd 3113 : data_o = 23'b 01001010100100110010100 ;
		12'd 3114 : data_o = 23'b 01001010011110111010111 ;
		12'd 3115 : data_o = 23'b 01001010011001000011100 ;
		12'd 3116 : data_o = 23'b 01001010010011001100010 ;
		12'd 3117 : data_o = 23'b 01001010001101010101001 ;
		12'd 3118 : data_o = 23'b 01001010000111011110010 ;
		12'd 3119 : data_o = 23'b 01001010000001100111011 ;
		12'd 3120 : data_o = 23'b 01001001111011110000110 ;
		12'd 3121 : data_o = 23'b 01001001110101111010010 ;
		12'd 3122 : data_o = 23'b 01001001110000000100000 ;
		12'd 3123 : data_o = 23'b 01001001101010001101110 ;
		12'd 3124 : data_o = 23'b 01001001100100010111110 ;
		12'd 3125 : data_o = 23'b 01001001011110100001111 ;
		12'd 3126 : data_o = 23'b 01001001011000101100010 ;
		12'd 3127 : data_o = 23'b 01001001010010110110101 ;
		12'd 3128 : data_o = 23'b 01001001001101000001010 ;
		12'd 3129 : data_o = 23'b 01001001000111001100000 ;
		12'd 3130 : data_o = 23'b 01001001000001010111000 ;
		12'd 3131 : data_o = 23'b 01001000111011100010000 ;
		12'd 3132 : data_o = 23'b 01001000110101101101010 ;
		12'd 3133 : data_o = 23'b 01001000101111111000101 ;
		12'd 3134 : data_o = 23'b 01001000101010000100001 ;
		12'd 3135 : data_o = 23'b 01001000100100001111111 ;
		12'd 3136 : data_o = 23'b 01001000011110011011110 ;
		12'd 3137 : data_o = 23'b 01001000011000100111110 ;
		12'd 3138 : data_o = 23'b 01001000010010110011111 ;
		12'd 3139 : data_o = 23'b 01001000001101000000001 ;
		12'd 3140 : data_o = 23'b 01001000000111001100101 ;
		12'd 3141 : data_o = 23'b 01001000000001011001010 ;
		12'd 3142 : data_o = 23'b 01000111111011100110000 ;
		12'd 3143 : data_o = 23'b 01000111110101110010111 ;
		12'd 3144 : data_o = 23'b 01000111110000000000000 ;
		12'd 3145 : data_o = 23'b 01000111101010001101010 ;
		12'd 3146 : data_o = 23'b 01000111100100011010101 ;
		12'd 3147 : data_o = 23'b 01000111011110101000001 ;
		12'd 3148 : data_o = 23'b 01000111011000110101111 ;
		12'd 3149 : data_o = 23'b 01000111010011000011101 ;
		12'd 3150 : data_o = 23'b 01000111001101010001101 ;
		12'd 3151 : data_o = 23'b 01000111000111011111111 ;
		12'd 3152 : data_o = 23'b 01000111000001101110001 ;
		12'd 3153 : data_o = 23'b 01000110111011111100101 ;
		12'd 3154 : data_o = 23'b 01000110110110001011010 ;
		12'd 3155 : data_o = 23'b 01000110110000011010000 ;
		12'd 3156 : data_o = 23'b 01000110101010101000111 ;
		12'd 3157 : data_o = 23'b 01000110100100111000000 ;
		12'd 3158 : data_o = 23'b 01000110011111000111001 ;
		12'd 3159 : data_o = 23'b 01000110011001010110100 ;
		12'd 3160 : data_o = 23'b 01000110010011100110001 ;
		12'd 3161 : data_o = 23'b 01000110001101110101110 ;
		12'd 3162 : data_o = 23'b 01000110001000000101101 ;
		12'd 3163 : data_o = 23'b 01000110000010010101100 ;
		12'd 3164 : data_o = 23'b 01000101111100100101110 ;
		12'd 3165 : data_o = 23'b 01000101110110110110000 ;
		12'd 3166 : data_o = 23'b 01000101110001000110011 ;
		12'd 3167 : data_o = 23'b 01000101101011010111000 ;
		12'd 3168 : data_o = 23'b 01000101100101100111110 ;
		12'd 3169 : data_o = 23'b 01000101011111111000101 ;
		12'd 3170 : data_o = 23'b 01000101011010001001101 ;
		12'd 3171 : data_o = 23'b 01000101010100011010111 ;
		12'd 3172 : data_o = 23'b 01000101001110101100010 ;
		12'd 3173 : data_o = 23'b 01000101001000111101110 ;
		12'd 3174 : data_o = 23'b 01000101000011001111011 ;
		12'd 3175 : data_o = 23'b 01000100111101100001001 ;
		12'd 3176 : data_o = 23'b 01000100110111110011001 ;
		12'd 3177 : data_o = 23'b 01000100110010000101010 ;
		12'd 3178 : data_o = 23'b 01000100101100010111100 ;
		12'd 3179 : data_o = 23'b 01000100100110101001111 ;
		12'd 3180 : data_o = 23'b 01000100100000111100100 ;
		12'd 3181 : data_o = 23'b 01000100011011001111001 ;
		12'd 3182 : data_o = 23'b 01000100010101100010000 ;
		12'd 3183 : data_o = 23'b 01000100001111110101000 ;
		12'd 3184 : data_o = 23'b 01000100001010001000001 ;
		12'd 3185 : data_o = 23'b 01000100000100011011100 ;
		12'd 3186 : data_o = 23'b 01000011111110101111000 ;
		12'd 3187 : data_o = 23'b 01000011111001000010100 ;
		12'd 3188 : data_o = 23'b 01000011110011010110010 ;
		12'd 3189 : data_o = 23'b 01000011101101101010010 ;
		12'd 3190 : data_o = 23'b 01000011100111111110010 ;
		12'd 3191 : data_o = 23'b 01000011100010010010100 ;
		12'd 3192 : data_o = 23'b 01000011011100100110111 ;
		12'd 3193 : data_o = 23'b 01000011010110111011011 ;
		12'd 3194 : data_o = 23'b 01000011010001010000000 ;
		12'd 3195 : data_o = 23'b 01000011001011100100111 ;
		12'd 3196 : data_o = 23'b 01000011000101111001110 ;
		12'd 3197 : data_o = 23'b 01000011000000001110111 ;
		12'd 3198 : data_o = 23'b 01000010111010100100001 ;
		12'd 3199 : data_o = 23'b 01000010110100111001100 ;
		12'd 3200 : data_o = 23'b 01000010101111001111001 ;
		12'd 3201 : data_o = 23'b 01000010101001100100110 ;
		12'd 3202 : data_o = 23'b 01000010100011111010101 ;
		12'd 3203 : data_o = 23'b 01000010011110010000101 ;
		12'd 3204 : data_o = 23'b 01000010011000100110110 ;
		12'd 3205 : data_o = 23'b 01000010010010111101001 ;
		12'd 3206 : data_o = 23'b 01000010001101010011100 ;
		12'd 3207 : data_o = 23'b 01000010000111101010001 ;
		12'd 3208 : data_o = 23'b 01000010000010000000111 ;
		12'd 3209 : data_o = 23'b 01000001111100010111110 ;
		12'd 3210 : data_o = 23'b 01000001110110101110110 ;
		12'd 3211 : data_o = 23'b 01000001110001000110000 ;
		12'd 3212 : data_o = 23'b 01000001101011011101011 ;
		12'd 3213 : data_o = 23'b 01000001100101110100110 ;
		12'd 3214 : data_o = 23'b 01000001100000001100011 ;
		12'd 3215 : data_o = 23'b 01000001011010100100010 ;
		12'd 3216 : data_o = 23'b 01000001010100111100001 ;
		12'd 3217 : data_o = 23'b 01000001001111010100010 ;
		12'd 3218 : data_o = 23'b 01000001001001101100100 ;
		12'd 3219 : data_o = 23'b 01000001000100000100110 ;
		12'd 3220 : data_o = 23'b 01000000111110011101011 ;
		12'd 3221 : data_o = 23'b 01000000111000110110000 ;
		12'd 3222 : data_o = 23'b 01000000110011001110110 ;
		12'd 3223 : data_o = 23'b 01000000101101100111110 ;
		12'd 3224 : data_o = 23'b 01000000101000000000111 ;
		12'd 3225 : data_o = 23'b 01000000100010011010001 ;
		12'd 3226 : data_o = 23'b 01000000011100110011100 ;
		12'd 3227 : data_o = 23'b 01000000010111001101001 ;
		12'd 3228 : data_o = 23'b 01000000010001100110110 ;
		12'd 3229 : data_o = 23'b 01000000001100000000101 ;
		12'd 3230 : data_o = 23'b 01000000000110011010101 ;
		12'd 3231 : data_o = 23'b 01000000000000110100110 ;
		12'd 3232 : data_o = 23'b 00111111111011001111000 ;
		12'd 3233 : data_o = 23'b 00111111110101101001011 ;
		12'd 3234 : data_o = 23'b 00111111110000000100000 ;
		12'd 3235 : data_o = 23'b 00111111101010011110110 ;
		12'd 3236 : data_o = 23'b 00111111100100111001101 ;
		12'd 3237 : data_o = 23'b 00111111011111010100101 ;
		12'd 3238 : data_o = 23'b 00111111011001101111110 ;
		12'd 3239 : data_o = 23'b 00111111010100001011001 ;
		12'd 3240 : data_o = 23'b 00111111001110100110100 ;
		12'd 3241 : data_o = 23'b 00111111001001000010001 ;
		12'd 3242 : data_o = 23'b 00111111000011011101111 ;
		12'd 3243 : data_o = 23'b 00111110111101111001110 ;
		12'd 3244 : data_o = 23'b 00111110111000010101110 ;
		12'd 3245 : data_o = 23'b 00111110110010110010000 ;
		12'd 3246 : data_o = 23'b 00111110101101001110010 ;
		12'd 3247 : data_o = 23'b 00111110100111101010110 ;
		12'd 3248 : data_o = 23'b 00111110100010000111011 ;
		12'd 3249 : data_o = 23'b 00111110011100100100001 ;
		12'd 3250 : data_o = 23'b 00111110010111000001000 ;
		12'd 3251 : data_o = 23'b 00111110010001011110001 ;
		12'd 3252 : data_o = 23'b 00111110001011111011010 ;
		12'd 3253 : data_o = 23'b 00111110000110011000101 ;
		12'd 3254 : data_o = 23'b 00111110000000110110001 ;
		12'd 3255 : data_o = 23'b 00111101111011010011110 ;
		12'd 3256 : data_o = 23'b 00111101110101110001100 ;
		12'd 3257 : data_o = 23'b 00111101110000001111011 ;
		12'd 3258 : data_o = 23'b 00111101101010101101100 ;
		12'd 3259 : data_o = 23'b 00111101100101001011101 ;
		12'd 3260 : data_o = 23'b 00111101011111101010000 ;
		12'd 3261 : data_o = 23'b 00111101011010001000100 ;
		12'd 3262 : data_o = 23'b 00111101010100100111001 ;
		12'd 3263 : data_o = 23'b 00111101001111000110000 ;
		12'd 3264 : data_o = 23'b 00111101001001100100111 ;
		12'd 3265 : data_o = 23'b 00111101000100000011111 ;
		12'd 3266 : data_o = 23'b 00111100111110100011001 ;
		12'd 3267 : data_o = 23'b 00111100111001000010100 ;
		12'd 3268 : data_o = 23'b 00111100110011100010000 ;
		12'd 3269 : data_o = 23'b 00111100101110000001101 ;
		12'd 3270 : data_o = 23'b 00111100101000100001100 ;
		12'd 3271 : data_o = 23'b 00111100100011000001011 ;
		12'd 3272 : data_o = 23'b 00111100011101100001100 ;
		12'd 3273 : data_o = 23'b 00111100011000000001101 ;
		12'd 3274 : data_o = 23'b 00111100010010100010000 ;
		12'd 3275 : data_o = 23'b 00111100001101000010100 ;
		12'd 3276 : data_o = 23'b 00111100000111100011010 ;
		12'd 3277 : data_o = 23'b 00111100000010000100000 ;
		12'd 3278 : data_o = 23'b 00111011111100100100111 ;
		12'd 3279 : data_o = 23'b 00111011110111000110000 ;
		12'd 3280 : data_o = 23'b 00111011110001100111010 ;
		12'd 3281 : data_o = 23'b 00111011101100001000101 ;
		12'd 3282 : data_o = 23'b 00111011100110101010001 ;
		12'd 3283 : data_o = 23'b 00111011100001001011110 ;
		12'd 3284 : data_o = 23'b 00111011011011101101100 ;
		12'd 3285 : data_o = 23'b 00111011010110001111100 ;
		12'd 3286 : data_o = 23'b 00111011010000110001100 ;
		12'd 3287 : data_o = 23'b 00111011001011010011110 ;
		12'd 3288 : data_o = 23'b 00111011000101110110001 ;
		12'd 3289 : data_o = 23'b 00111011000000011000101 ;
		12'd 3290 : data_o = 23'b 00111010111010111011010 ;
		12'd 3291 : data_o = 23'b 00111010110101011110000 ;
		12'd 3292 : data_o = 23'b 00111010110000000001000 ;
		12'd 3293 : data_o = 23'b 00111010101010100100000 ;
		12'd 3294 : data_o = 23'b 00111010100101000111010 ;
		12'd 3295 : data_o = 23'b 00111010011111101010101 ;
		12'd 3296 : data_o = 23'b 00111010011010001110001 ;
		12'd 3297 : data_o = 23'b 00111010010100110001110 ;
		12'd 3298 : data_o = 23'b 00111010001111010101100 ;
		12'd 3299 : data_o = 23'b 00111010001001111001011 ;
		12'd 3300 : data_o = 23'b 00111010000100011101100 ;
		12'd 3301 : data_o = 23'b 00111001111111000001101 ;
		12'd 3302 : data_o = 23'b 00111001111001100110000 ;
		12'd 3303 : data_o = 23'b 00111001110100001010100 ;
		12'd 3304 : data_o = 23'b 00111001101110101111001 ;
		12'd 3305 : data_o = 23'b 00111001101001010011111 ;
		12'd 3306 : data_o = 23'b 00111001100011111000110 ;
		12'd 3307 : data_o = 23'b 00111001011110011101110 ;
		12'd 3308 : data_o = 23'b 00111001011001000011000 ;
		12'd 3309 : data_o = 23'b 00111001010011101000010 ;
		12'd 3310 : data_o = 23'b 00111001001110001101110 ;
		12'd 3311 : data_o = 23'b 00111001001000110011011 ;
		12'd 3312 : data_o = 23'b 00111001000011011001001 ;
		12'd 3313 : data_o = 23'b 00111000111101111111000 ;
		12'd 3314 : data_o = 23'b 00111000111000100101000 ;
		12'd 3315 : data_o = 23'b 00111000110011001011010 ;
		12'd 3316 : data_o = 23'b 00111000101101110001100 ;
		12'd 3317 : data_o = 23'b 00111000101000011000000 ;
		12'd 3318 : data_o = 23'b 00111000100010111110100 ;
		12'd 3319 : data_o = 23'b 00111000011101100101010 ;
		12'd 3320 : data_o = 23'b 00111000011000001100001 ;
		12'd 3321 : data_o = 23'b 00111000010010110011001 ;
		12'd 3322 : data_o = 23'b 00111000001101011010010 ;
		12'd 3323 : data_o = 23'b 00111000001000000001101 ;
		12'd 3324 : data_o = 23'b 00111000000010101001000 ;
		12'd 3325 : data_o = 23'b 00110111111101010000100 ;
		12'd 3326 : data_o = 23'b 00110111110111111000010 ;
		12'd 3327 : data_o = 23'b 00110111110010100000001 ;
		12'd 3328 : data_o = 23'b 00110111101101001000001 ;
		12'd 3329 : data_o = 23'b 00110111100111110000010 ;
		12'd 3330 : data_o = 23'b 00110111100010011000100 ;
		12'd 3331 : data_o = 23'b 00110111011101000000111 ;
		12'd 3332 : data_o = 23'b 00110111010111101001011 ;
		12'd 3333 : data_o = 23'b 00110111010010010010001 ;
		12'd 3334 : data_o = 23'b 00110111001100111010111 ;
		12'd 3335 : data_o = 23'b 00110111000111100011111 ;
		12'd 3336 : data_o = 23'b 00110111000010001100111 ;
		12'd 3337 : data_o = 23'b 00110110111100110110001 ;
		12'd 3338 : data_o = 23'b 00110110110111011111100 ;
		12'd 3339 : data_o = 23'b 00110110110010001001000 ;
		12'd 3340 : data_o = 23'b 00110110101100110010101 ;
		12'd 3341 : data_o = 23'b 00110110100111011100100 ;
		12'd 3342 : data_o = 23'b 00110110100010000110011 ;
		12'd 3343 : data_o = 23'b 00110110011100110000011 ;
		12'd 3344 : data_o = 23'b 00110110010111011010101 ;
		12'd 3345 : data_o = 23'b 00110110010010000101000 ;
		12'd 3346 : data_o = 23'b 00110110001100101111011 ;
		12'd 3347 : data_o = 23'b 00110110000111011010000 ;
		12'd 3348 : data_o = 23'b 00110110000010000100110 ;
		12'd 3349 : data_o = 23'b 00110101111100101111101 ;
		12'd 3350 : data_o = 23'b 00110101110111011010101 ;
		12'd 3351 : data_o = 23'b 00110101110010000101111 ;
		12'd 3352 : data_o = 23'b 00110101101100110001001 ;
		12'd 3353 : data_o = 23'b 00110101100111011100100 ;
		12'd 3354 : data_o = 23'b 00110101100010001000001 ;
		12'd 3355 : data_o = 23'b 00110101011100110011111 ;
		12'd 3356 : data_o = 23'b 00110101010111011111101 ;
		12'd 3357 : data_o = 23'b 00110101010010001011101 ;
		12'd 3358 : data_o = 23'b 00110101001100110111110 ;
		12'd 3359 : data_o = 23'b 00110101000111100100000 ;
		12'd 3360 : data_o = 23'b 00110101000010010000011 ;
		12'd 3361 : data_o = 23'b 00110100111100111101000 ;
		12'd 3362 : data_o = 23'b 00110100110111101001101 ;
		12'd 3363 : data_o = 23'b 00110100110010010110011 ;
		12'd 3364 : data_o = 23'b 00110100101101000011011 ;
		12'd 3365 : data_o = 23'b 00110100100111110000011 ;
		12'd 3366 : data_o = 23'b 00110100100010011101101 ;
		12'd 3367 : data_o = 23'b 00110100011101001011000 ;
		12'd 3368 : data_o = 23'b 00110100010111111000100 ;
		12'd 3369 : data_o = 23'b 00110100010010100110001 ;
		12'd 3370 : data_o = 23'b 00110100001101010011111 ;
		12'd 3371 : data_o = 23'b 00110100001000000001110 ;
		12'd 3372 : data_o = 23'b 00110100000010101111110 ;
		12'd 3373 : data_o = 23'b 00110011111101011101111 ;
		12'd 3374 : data_o = 23'b 00110011111000001100010 ;
		12'd 3375 : data_o = 23'b 00110011110010111010101 ;
		12'd 3376 : data_o = 23'b 00110011101101101001010 ;
		12'd 3377 : data_o = 23'b 00110011101000010111111 ;
		12'd 3378 : data_o = 23'b 00110011100011000110110 ;
		12'd 3379 : data_o = 23'b 00110011011101110101110 ;
		12'd 3380 : data_o = 23'b 00110011011000100100111 ;
		12'd 3381 : data_o = 23'b 00110011010011010100001 ;
		12'd 3382 : data_o = 23'b 00110011001110000011100 ;
		12'd 3383 : data_o = 23'b 00110011001000110011000 ;
		12'd 3384 : data_o = 23'b 00110011000011100010101 ;
		12'd 3385 : data_o = 23'b 00110010111110010010011 ;
		12'd 3386 : data_o = 23'b 00110010111001000010011 ;
		12'd 3387 : data_o = 23'b 00110010110011110010011 ;
		12'd 3388 : data_o = 23'b 00110010101110100010101 ;
		12'd 3389 : data_o = 23'b 00110010101001010010111 ;
		12'd 3390 : data_o = 23'b 00110010100100000011011 ;
		12'd 3391 : data_o = 23'b 00110010011110110011111 ;
		12'd 3392 : data_o = 23'b 00110010011001100100101 ;
		12'd 3393 : data_o = 23'b 00110010010100010101100 ;
		12'd 3394 : data_o = 23'b 00110010001111000110100 ;
		12'd 3395 : data_o = 23'b 00110010001001110111101 ;
		12'd 3396 : data_o = 23'b 00110010000100101000111 ;
		12'd 3397 : data_o = 23'b 00110001111111011010010 ;
		12'd 3398 : data_o = 23'b 00110001111010001011111 ;
		12'd 3399 : data_o = 23'b 00110001110100111101100 ;
		12'd 3400 : data_o = 23'b 00110001101111101111010 ;
		12'd 3401 : data_o = 23'b 00110001101010100001010 ;
		12'd 3402 : data_o = 23'b 00110001100101010011010 ;
		12'd 3403 : data_o = 23'b 00110001100000000101100 ;
		12'd 3404 : data_o = 23'b 00110001011010110111111 ;
		12'd 3405 : data_o = 23'b 00110001010101101010010 ;
		12'd 3406 : data_o = 23'b 00110001010000011100111 ;
		12'd 3407 : data_o = 23'b 00110001001011001111101 ;
		12'd 3408 : data_o = 23'b 00110001000110000010100 ;
		12'd 3409 : data_o = 23'b 00110001000000110101100 ;
		12'd 3410 : data_o = 23'b 00110000111011101000101 ;
		12'd 3411 : data_o = 23'b 00110000110110011011111 ;
		12'd 3412 : data_o = 23'b 00110000110001001111010 ;
		12'd 3413 : data_o = 23'b 00110000101100000010111 ;
		12'd 3414 : data_o = 23'b 00110000100110110110100 ;
		12'd 3415 : data_o = 23'b 00110000100001101010010 ;
		12'd 3416 : data_o = 23'b 00110000011100011110010 ;
		12'd 3417 : data_o = 23'b 00110000010111010010010 ;
		12'd 3418 : data_o = 23'b 00110000010010000110100 ;
		12'd 3419 : data_o = 23'b 00110000001100111010110 ;
		12'd 3420 : data_o = 23'b 00110000000111101111010 ;
		12'd 3421 : data_o = 23'b 00110000000010100011111 ;
		12'd 3422 : data_o = 23'b 00101111111101011000101 ;
		12'd 3423 : data_o = 23'b 00101111111000001101100 ;
		12'd 3424 : data_o = 23'b 00101111110011000010011 ;
		12'd 3425 : data_o = 23'b 00101111101101110111100 ;
		12'd 3426 : data_o = 23'b 00101111101000101100110 ;
		12'd 3427 : data_o = 23'b 00101111100011100010001 ;
		12'd 3428 : data_o = 23'b 00101111011110010111110 ;
		12'd 3429 : data_o = 23'b 00101111011001001101011 ;
		12'd 3430 : data_o = 23'b 00101111010100000011001 ;
		12'd 3431 : data_o = 23'b 00101111001110111001000 ;
		12'd 3432 : data_o = 23'b 00101111001001101111001 ;
		12'd 3433 : data_o = 23'b 00101111000100100101010 ;
		12'd 3434 : data_o = 23'b 00101110111111011011101 ;
		12'd 3435 : data_o = 23'b 00101110111010010010000 ;
		12'd 3436 : data_o = 23'b 00101110110101001000101 ;
		12'd 3437 : data_o = 23'b 00101110101111111111010 ;
		12'd 3438 : data_o = 23'b 00101110101010110110001 ;
		12'd 3439 : data_o = 23'b 00101110100101101101000 ;
		12'd 3440 : data_o = 23'b 00101110100000100100001 ;
		12'd 3441 : data_o = 23'b 00101110011011011011011 ;
		12'd 3442 : data_o = 23'b 00101110010110010010110 ;
		12'd 3443 : data_o = 23'b 00101110010001001010010 ;
		12'd 3444 : data_o = 23'b 00101110001100000001111 ;
		12'd 3445 : data_o = 23'b 00101110000110111001101 ;
		12'd 3446 : data_o = 23'b 00101110000001110001100 ;
		12'd 3447 : data_o = 23'b 00101101111100101001100 ;
		12'd 3448 : data_o = 23'b 00101101110111100001101 ;
		12'd 3449 : data_o = 23'b 00101101110010011001111 ;
		12'd 3450 : data_o = 23'b 00101101101101010010010 ;
		12'd 3451 : data_o = 23'b 00101101101000001010110 ;
		12'd 3452 : data_o = 23'b 00101101100011000011100 ;
		12'd 3453 : data_o = 23'b 00101101011101111100010 ;
		12'd 3454 : data_o = 23'b 00101101011000110101001 ;
		12'd 3455 : data_o = 23'b 00101101010011101110010 ;
		12'd 3456 : data_o = 23'b 00101101001110100111011 ;
		12'd 3457 : data_o = 23'b 00101101001001100000110 ;
		12'd 3458 : data_o = 23'b 00101101000100011010001 ;
		12'd 3459 : data_o = 23'b 00101100111111010011110 ;
		12'd 3460 : data_o = 23'b 00101100111010001101011 ;
		12'd 3461 : data_o = 23'b 00101100110101000111010 ;
		12'd 3462 : data_o = 23'b 00101100110000000001010 ;
		12'd 3463 : data_o = 23'b 00101100101010111011010 ;
		12'd 3464 : data_o = 23'b 00101100100101110101100 ;
		12'd 3465 : data_o = 23'b 00101100100000101111111 ;
		12'd 3466 : data_o = 23'b 00101100011011101010010 ;
		12'd 3467 : data_o = 23'b 00101100010110100100111 ;
		12'd 3468 : data_o = 23'b 00101100010001011111101 ;
		12'd 3469 : data_o = 23'b 00101100001100011010100 ;
		12'd 3470 : data_o = 23'b 00101100000111010101100 ;
		12'd 3471 : data_o = 23'b 00101100000010010000101 ;
		12'd 3472 : data_o = 23'b 00101011111101001011111 ;
		12'd 3473 : data_o = 23'b 00101011111000000111010 ;
		12'd 3474 : data_o = 23'b 00101011110011000010110 ;
		12'd 3475 : data_o = 23'b 00101011101101111110011 ;
		12'd 3476 : data_o = 23'b 00101011101000111010001 ;
		12'd 3477 : data_o = 23'b 00101011100011110110000 ;
		12'd 3478 : data_o = 23'b 00101011011110110010000 ;
		12'd 3479 : data_o = 23'b 00101011011001101110010 ;
		12'd 3480 : data_o = 23'b 00101011010100101010100 ;
		12'd 3481 : data_o = 23'b 00101011001111100110111 ;
		12'd 3482 : data_o = 23'b 00101011001010100011011 ;
		12'd 3483 : data_o = 23'b 00101011000101100000001 ;
		12'd 3484 : data_o = 23'b 00101011000000011100111 ;
		12'd 3485 : data_o = 23'b 00101010111011011001110 ;
		12'd 3486 : data_o = 23'b 00101010110110010110110 ;
		12'd 3487 : data_o = 23'b 00101010110001010100000 ;
		12'd 3488 : data_o = 23'b 00101010101100010001010 ;
		12'd 3489 : data_o = 23'b 00101010100111001110110 ;
		12'd 3490 : data_o = 23'b 00101010100010001100010 ;
		12'd 3491 : data_o = 23'b 00101010011101001010000 ;
		12'd 3492 : data_o = 23'b 00101010011000000111110 ;
		12'd 3493 : data_o = 23'b 00101010010011000101101 ;
		12'd 3494 : data_o = 23'b 00101010001110000011110 ;
		12'd 3495 : data_o = 23'b 00101010001001000010000 ;
		12'd 3496 : data_o = 23'b 00101010000100000000010 ;
		12'd 3497 : data_o = 23'b 00101001111110111110110 ;
		12'd 3498 : data_o = 23'b 00101001111001111101010 ;
		12'd 3499 : data_o = 23'b 00101001110100111100000 ;
		12'd 3500 : data_o = 23'b 00101001101111111010110 ;
		12'd 3501 : data_o = 23'b 00101001101010111001110 ;
		12'd 3502 : data_o = 23'b 00101001100101111000111 ;
		12'd 3503 : data_o = 23'b 00101001100000111000000 ;
		12'd 3504 : data_o = 23'b 00101001011011110111011 ;
		12'd 3505 : data_o = 23'b 00101001010110110110111 ;
		12'd 3506 : data_o = 23'b 00101001010001110110011 ;
		12'd 3507 : data_o = 23'b 00101001001100110110001 ;
		12'd 3508 : data_o = 23'b 00101001000111110110000 ;
		12'd 3509 : data_o = 23'b 00101001000010110101111 ;
		12'd 3510 : data_o = 23'b 00101000111101110110000 ;
		12'd 3511 : data_o = 23'b 00101000111000110110010 ;
		12'd 3512 : data_o = 23'b 00101000110011110110101 ;
		12'd 3513 : data_o = 23'b 00101000101110110111000 ;
		12'd 3514 : data_o = 23'b 00101000101001110111101 ;
		12'd 3515 : data_o = 23'b 00101000100100111000011 ;
		12'd 3516 : data_o = 23'b 00101000011111111001010 ;
		12'd 3517 : data_o = 23'b 00101000011010111010001 ;
		12'd 3518 : data_o = 23'b 00101000010101111011010 ;
		12'd 3519 : data_o = 23'b 00101000010000111100100 ;
		12'd 3520 : data_o = 23'b 00101000001011111101111 ;
		12'd 3521 : data_o = 23'b 00101000000110111111011 ;
		12'd 3522 : data_o = 23'b 00101000000010000000111 ;
		12'd 3523 : data_o = 23'b 00100111111101000010101 ;
		12'd 3524 : data_o = 23'b 00100111111000000100100 ;
		12'd 3525 : data_o = 23'b 00100111110011000110100 ;
		12'd 3526 : data_o = 23'b 00100111101110001000101 ;
		12'd 3527 : data_o = 23'b 00100111101001001010111 ;
		12'd 3528 : data_o = 23'b 00100111100100001101001 ;
		12'd 3529 : data_o = 23'b 00100111011111001111101 ;
		12'd 3530 : data_o = 23'b 00100111011010010010010 ;
		12'd 3531 : data_o = 23'b 00100111010101010101000 ;
		12'd 3532 : data_o = 23'b 00100111010000010111111 ;
		12'd 3533 : data_o = 23'b 00100111001011011010110 ;
		12'd 3534 : data_o = 23'b 00100111000110011101111 ;
		12'd 3535 : data_o = 23'b 00100111000001100001001 ;
		12'd 3536 : data_o = 23'b 00100110111100100100100 ;
		12'd 3537 : data_o = 23'b 00100110110111101000000 ;
		12'd 3538 : data_o = 23'b 00100110110010101011100 ;
		12'd 3539 : data_o = 23'b 00100110101101101111010 ;
		12'd 3540 : data_o = 23'b 00100110101000110011001 ;
		12'd 3541 : data_o = 23'b 00100110100011110111001 ;
		12'd 3542 : data_o = 23'b 00100110011110111011001 ;
		12'd 3543 : data_o = 23'b 00100110011001111111011 ;
		12'd 3544 : data_o = 23'b 00100110010101000011110 ;
		12'd 3545 : data_o = 23'b 00100110010000001000010 ;
		12'd 3546 : data_o = 23'b 00100110001011001100110 ;
		12'd 3547 : data_o = 23'b 00100110000110010001100 ;
		12'd 3548 : data_o = 23'b 00100110000001010110011 ;
		12'd 3549 : data_o = 23'b 00100101111100011011011 ;
		12'd 3550 : data_o = 23'b 00100101110111100000011 ;
		12'd 3551 : data_o = 23'b 00100101110010100101101 ;
		12'd 3552 : data_o = 23'b 00100101101101101011000 ;
		12'd 3553 : data_o = 23'b 00100101101000110000011 ;
		12'd 3554 : data_o = 23'b 00100101100011110110000 ;
		12'd 3555 : data_o = 23'b 00100101011110111011101 ;
		12'd 3556 : data_o = 23'b 00100101011010000001100 ;
		12'd 3557 : data_o = 23'b 00100101010101000111100 ;
		12'd 3558 : data_o = 23'b 00100101010000001101100 ;
		12'd 3559 : data_o = 23'b 00100101001011010011110 ;
		12'd 3560 : data_o = 23'b 00100101000110011010000 ;
		12'd 3561 : data_o = 23'b 00100101000001100000100 ;
		12'd 3562 : data_o = 23'b 00100100111100100111000 ;
		12'd 3563 : data_o = 23'b 00100100110111101101110 ;
		12'd 3564 : data_o = 23'b 00100100110010110100100 ;
		12'd 3565 : data_o = 23'b 00100100101101111011100 ;
		12'd 3566 : data_o = 23'b 00100100101001000010100 ;
		12'd 3567 : data_o = 23'b 00100100100100001001110 ;
		12'd 3568 : data_o = 23'b 00100100011111010001000 ;
		12'd 3569 : data_o = 23'b 00100100011010011000011 ;
		12'd 3570 : data_o = 23'b 00100100010101100000000 ;
		12'd 3571 : data_o = 23'b 00100100010000100111101 ;
		12'd 3572 : data_o = 23'b 00100100001011101111011 ;
		12'd 3573 : data_o = 23'b 00100100000110110111011 ;
		12'd 3574 : data_o = 23'b 00100100000001111111011 ;
		12'd 3575 : data_o = 23'b 00100011111101000111100 ;
		12'd 3576 : data_o = 23'b 00100011111000001111110 ;
		12'd 3577 : data_o = 23'b 00100011110011011000010 ;
		12'd 3578 : data_o = 23'b 00100011101110100000110 ;
		12'd 3579 : data_o = 23'b 00100011101001101001011 ;
		12'd 3580 : data_o = 23'b 00100011100100110010001 ;
		12'd 3581 : data_o = 23'b 00100011011111111011000 ;
		12'd 3582 : data_o = 23'b 00100011011011000100000 ;
		12'd 3583 : data_o = 23'b 00100011010110001101001 ;
		12'd 3584 : data_o = 23'b 00100011010001010110011 ;
		12'd 3585 : data_o = 23'b 00100011001100011111110 ;
		12'd 3586 : data_o = 23'b 00100011000111101001010 ;
		12'd 3587 : data_o = 23'b 00100011000010110010111 ;
		12'd 3588 : data_o = 23'b 00100010111101111100101 ;
		12'd 3589 : data_o = 23'b 00100010111001000110100 ;
		12'd 3590 : data_o = 23'b 00100010110100010000100 ;
		12'd 3591 : data_o = 23'b 00100010101111011010100 ;
		12'd 3592 : data_o = 23'b 00100010101010100100110 ;
		12'd 3593 : data_o = 23'b 00100010100101101111001 ;
		12'd 3594 : data_o = 23'b 00100010100000111001101 ;
		12'd 3595 : data_o = 23'b 00100010011100000100001 ;
		12'd 3596 : data_o = 23'b 00100010010111001110111 ;
		12'd 3597 : data_o = 23'b 00100010010010011001101 ;
		12'd 3598 : data_o = 23'b 00100010001101100100101 ;
		12'd 3599 : data_o = 23'b 00100010001000101111110 ;
		12'd 3600 : data_o = 23'b 00100010000011111010111 ;
		12'd 3601 : data_o = 23'b 00100001111111000110001 ;
		12'd 3602 : data_o = 23'b 00100001111010010001101 ;
		12'd 3603 : data_o = 23'b 00100001110101011101001 ;
		12'd 3604 : data_o = 23'b 00100001110000101000111 ;
		12'd 3605 : data_o = 23'b 00100001101011110100101 ;
		12'd 3606 : data_o = 23'b 00100001100111000000100 ;
		12'd 3607 : data_o = 23'b 00100001100010001100100 ;
		12'd 3608 : data_o = 23'b 00100001011101011000101 ;
		12'd 3609 : data_o = 23'b 00100001011000100101000 ;
		12'd 3610 : data_o = 23'b 00100001010011110001011 ;
		12'd 3611 : data_o = 23'b 00100001001110111101111 ;
		12'd 3612 : data_o = 23'b 00100001001010001010100 ;
		12'd 3613 : data_o = 23'b 00100001000101010111010 ;
		12'd 3614 : data_o = 23'b 00100001000000100100001 ;
		12'd 3615 : data_o = 23'b 00100000111011110001000 ;
		12'd 3616 : data_o = 23'b 00100000110110111110001 ;
		12'd 3617 : data_o = 23'b 00100000110010001011011 ;
		12'd 3618 : data_o = 23'b 00100000101101011000110 ;
		12'd 3619 : data_o = 23'b 00100000101000100110001 ;
		12'd 3620 : data_o = 23'b 00100000100011110011110 ;
		12'd 3621 : data_o = 23'b 00100000011111000001100 ;
		12'd 3622 : data_o = 23'b 00100000011010001111010 ;
		12'd 3623 : data_o = 23'b 00100000010101011101010 ;
		12'd 3624 : data_o = 23'b 00100000010000101011010 ;
		12'd 3625 : data_o = 23'b 00100000001011111001011 ;
		12'd 3626 : data_o = 23'b 00100000000111000111110 ;
		12'd 3627 : data_o = 23'b 00100000000010010110001 ;
		12'd 3628 : data_o = 23'b 00011111111101100100101 ;
		12'd 3629 : data_o = 23'b 00011111111000110011011 ;
		12'd 3630 : data_o = 23'b 00011111110100000010001 ;
		12'd 3631 : data_o = 23'b 00011111101111010001000 ;
		12'd 3632 : data_o = 23'b 00011111101010100000000 ;
		12'd 3633 : data_o = 23'b 00011111100101101111001 ;
		12'd 3634 : data_o = 23'b 00011111100000111110011 ;
		12'd 3635 : data_o = 23'b 00011111011100001101110 ;
		12'd 3636 : data_o = 23'b 00011111010111011101001 ;
		12'd 3637 : data_o = 23'b 00011111010010101100110 ;
		12'd 3638 : data_o = 23'b 00011111001101111100100 ;
		12'd 3639 : data_o = 23'b 00011111001001001100011 ;
		12'd 3640 : data_o = 23'b 00011111000100011100010 ;
		12'd 3641 : data_o = 23'b 00011110111111101100011 ;
		12'd 3642 : data_o = 23'b 00011110111010111100100 ;
		12'd 3643 : data_o = 23'b 00011110110110001100111 ;
		12'd 3644 : data_o = 23'b 00011110110001011101010 ;
		12'd 3645 : data_o = 23'b 00011110101100101101110 ;
		12'd 3646 : data_o = 23'b 00011110100111111110100 ;
		12'd 3647 : data_o = 23'b 00011110100011001111010 ;
		12'd 3648 : data_o = 23'b 00011110011110100000001 ;
		12'd 3649 : data_o = 23'b 00011110011001110001001 ;
		12'd 3650 : data_o = 23'b 00011110010101000010010 ;
		12'd 3651 : data_o = 23'b 00011110010000010011100 ;
		12'd 3652 : data_o = 23'b 00011110001011100100111 ;
		12'd 3653 : data_o = 23'b 00011110000110110110011 ;
		12'd 3654 : data_o = 23'b 00011110000010000111111 ;
		12'd 3655 : data_o = 23'b 00011101111101011001101 ;
		12'd 3656 : data_o = 23'b 00011101111000101011100 ;
		12'd 3657 : data_o = 23'b 00011101110011111101011 ;
		12'd 3658 : data_o = 23'b 00011101101111001111100 ;
		12'd 3659 : data_o = 23'b 00011101101010100001101 ;
		12'd 3660 : data_o = 23'b 00011101100101110100000 ;
		12'd 3661 : data_o = 23'b 00011101100001000110011 ;
		12'd 3662 : data_o = 23'b 00011101011100011000111 ;
		12'd 3663 : data_o = 23'b 00011101010111101011100 ;
		12'd 3664 : data_o = 23'b 00011101010010111110010 ;
		12'd 3665 : data_o = 23'b 00011101001110010001010 ;
		12'd 3666 : data_o = 23'b 00011101001001100100001 ;
		12'd 3667 : data_o = 23'b 00011101000100110111010 ;
		12'd 3668 : data_o = 23'b 00011101000000001010100 ;
		12'd 3669 : data_o = 23'b 00011100111011011101111 ;
		12'd 3670 : data_o = 23'b 00011100110110110001011 ;
		12'd 3671 : data_o = 23'b 00011100110010000100111 ;
		12'd 3672 : data_o = 23'b 00011100101101011000101 ;
		12'd 3673 : data_o = 23'b 00011100101000101100011 ;
		12'd 3674 : data_o = 23'b 00011100100100000000011 ;
		12'd 3675 : data_o = 23'b 00011100011111010100011 ;
		12'd 3676 : data_o = 23'b 00011100011010101000100 ;
		12'd 3677 : data_o = 23'b 00011100010101111100110 ;
		12'd 3678 : data_o = 23'b 00011100010001010001010 ;
		12'd 3679 : data_o = 23'b 00011100001100100101110 ;
		12'd 3680 : data_o = 23'b 00011100000111111010010 ;
		12'd 3681 : data_o = 23'b 00011100000011001111000 ;
		12'd 3682 : data_o = 23'b 00011011111110100011111 ;
		12'd 3683 : data_o = 23'b 00011011111001111000111 ;
		12'd 3684 : data_o = 23'b 00011011110101001110000 ;
		12'd 3685 : data_o = 23'b 00011011110000100011001 ;
		12'd 3686 : data_o = 23'b 00011011101011111000100 ;
		12'd 3687 : data_o = 23'b 00011011100111001101111 ;
		12'd 3688 : data_o = 23'b 00011011100010100011011 ;
		12'd 3689 : data_o = 23'b 00011011011101111001001 ;
		12'd 3690 : data_o = 23'b 00011011011001001110111 ;
		12'd 3691 : data_o = 23'b 00011011010100100100110 ;
		12'd 3692 : data_o = 23'b 00011011001111111010110 ;
		12'd 3693 : data_o = 23'b 00011011001011010000111 ;
		12'd 3694 : data_o = 23'b 00011011000110100111001 ;
		12'd 3695 : data_o = 23'b 00011011000001111101011 ;
		12'd 3696 : data_o = 23'b 00011010111101010011111 ;
		12'd 3697 : data_o = 23'b 00011010111000101010100 ;
		12'd 3698 : data_o = 23'b 00011010110100000001001 ;
		12'd 3699 : data_o = 23'b 00011010101111010111111 ;
		12'd 3700 : data_o = 23'b 00011010101010101110111 ;
		12'd 3701 : data_o = 23'b 00011010100110000101111 ;
		12'd 3702 : data_o = 23'b 00011010100001011101000 ;
		12'd 3703 : data_o = 23'b 00011010011100110100010 ;
		12'd 3704 : data_o = 23'b 00011010011000001011101 ;
		12'd 3705 : data_o = 23'b 00011010010011100011001 ;
		12'd 3706 : data_o = 23'b 00011010001110111010110 ;
		12'd 3707 : data_o = 23'b 00011010001010010010100 ;
		12'd 3708 : data_o = 23'b 00011010000101101010010 ;
		12'd 3709 : data_o = 23'b 00011010000001000010010 ;
		12'd 3710 : data_o = 23'b 00011001111100011010010 ;
		12'd 3711 : data_o = 23'b 00011001110111110010100 ;
		12'd 3712 : data_o = 23'b 00011001110011001010110 ;
		12'd 3713 : data_o = 23'b 00011001101110100011001 ;
		12'd 3714 : data_o = 23'b 00011001101001111011101 ;
		12'd 3715 : data_o = 23'b 00011001100101010100010 ;
		12'd 3716 : data_o = 23'b 00011001100000101101000 ;
		12'd 3717 : data_o = 23'b 00011001011100000101111 ;
		12'd 3718 : data_o = 23'b 00011001010111011110111 ;
		12'd 3719 : data_o = 23'b 00011001010010110111111 ;
		12'd 3720 : data_o = 23'b 00011001001110010001001 ;
		12'd 3721 : data_o = 23'b 00011001001001101010011 ;
		12'd 3722 : data_o = 23'b 00011001000101000011111 ;
		12'd 3723 : data_o = 23'b 00011001000000011101011 ;
		12'd 3724 : data_o = 23'b 00011000111011110111000 ;
		12'd 3725 : data_o = 23'b 00011000110111010000110 ;
		12'd 3726 : data_o = 23'b 00011000110010101010101 ;
		12'd 3727 : data_o = 23'b 00011000101110000100101 ;
		12'd 3728 : data_o = 23'b 00011000101001011110110 ;
		12'd 3729 : data_o = 23'b 00011000100100111000111 ;
		12'd 3730 : data_o = 23'b 00011000100000010011010 ;
		12'd 3731 : data_o = 23'b 00011000011011101101101 ;
		12'd 3732 : data_o = 23'b 00011000010111001000010 ;
		12'd 3733 : data_o = 23'b 00011000010010100010111 ;
		12'd 3734 : data_o = 23'b 00011000001101111101101 ;
		12'd 3735 : data_o = 23'b 00011000001001011000100 ;
		12'd 3736 : data_o = 23'b 00011000000100110011100 ;
		12'd 3737 : data_o = 23'b 00011000000000001110101 ;
		12'd 3738 : data_o = 23'b 00010111111011101001111 ;
		12'd 3739 : data_o = 23'b 00010111110111000101010 ;
		12'd 3740 : data_o = 23'b 00010111110010100000101 ;
		12'd 3741 : data_o = 23'b 00010111101101111100010 ;
		12'd 3742 : data_o = 23'b 00010111101001010111111 ;
		12'd 3743 : data_o = 23'b 00010111100100110011101 ;
		12'd 3744 : data_o = 23'b 00010111100000001111100 ;
		12'd 3745 : data_o = 23'b 00010111011011101011100 ;
		12'd 3746 : data_o = 23'b 00010111010111000111101 ;
		12'd 3747 : data_o = 23'b 00010111010010100011111 ;
		12'd 3748 : data_o = 23'b 00010111001110000000010 ;
		12'd 3749 : data_o = 23'b 00010111001001011100101 ;
		12'd 3750 : data_o = 23'b 00010111000100111001010 ;
		12'd 3751 : data_o = 23'b 00010111000000010101111 ;
		12'd 3752 : data_o = 23'b 00010110111011110010101 ;
		12'd 3753 : data_o = 23'b 00010110110111001111101 ;
		12'd 3754 : data_o = 23'b 00010110110010101100101 ;
		12'd 3755 : data_o = 23'b 00010110101110001001110 ;
		12'd 3756 : data_o = 23'b 00010110101001100110111 ;
		12'd 3757 : data_o = 23'b 00010110100101000100010 ;
		12'd 3758 : data_o = 23'b 00010110100000100001110 ;
		12'd 3759 : data_o = 23'b 00010110011011111111010 ;
		12'd 3760 : data_o = 23'b 00010110010111011101000 ;
		12'd 3761 : data_o = 23'b 00010110010010111010110 ;
		12'd 3762 : data_o = 23'b 00010110001110011000101 ;
		12'd 3763 : data_o = 23'b 00010110001001110110101 ;
		12'd 3764 : data_o = 23'b 00010110000101010100110 ;
		12'd 3765 : data_o = 23'b 00010110000000110011000 ;
		12'd 3766 : data_o = 23'b 00010101111100010001010 ;
		12'd 3767 : data_o = 23'b 00010101110111101111110 ;
		12'd 3768 : data_o = 23'b 00010101110011001110011 ;
		12'd 3769 : data_o = 23'b 00010101101110101101000 ;
		12'd 3770 : data_o = 23'b 00010101101010001011110 ;
		12'd 3771 : data_o = 23'b 00010101100101101010101 ;
		12'd 3772 : data_o = 23'b 00010101100001001001101 ;
		12'd 3773 : data_o = 23'b 00010101011100101000110 ;
		12'd 3774 : data_o = 23'b 00010101011000001000000 ;
		12'd 3775 : data_o = 23'b 00010101010011100111010 ;
		12'd 3776 : data_o = 23'b 00010101001111000110110 ;
		12'd 3777 : data_o = 23'b 00010101001010100110010 ;
		12'd 3778 : data_o = 23'b 00010101000110000110000 ;
		12'd 3779 : data_o = 23'b 00010101000001100101110 ;
		12'd 3780 : data_o = 23'b 00010100111101000101101 ;
		12'd 3781 : data_o = 23'b 00010100111000100101101 ;
		12'd 3782 : data_o = 23'b 00010100110100000101101 ;
		12'd 3783 : data_o = 23'b 00010100101111100101111 ;
		12'd 3784 : data_o = 23'b 00010100101011000110010 ;
		12'd 3785 : data_o = 23'b 00010100100110100110101 ;
		12'd 3786 : data_o = 23'b 00010100100010000111001 ;
		12'd 3787 : data_o = 23'b 00010100011101100111111 ;
		12'd 3788 : data_o = 23'b 00010100011001001000101 ;
		12'd 3789 : data_o = 23'b 00010100010100101001100 ;
		12'd 3790 : data_o = 23'b 00010100010000001010011 ;
		12'd 3791 : data_o = 23'b 00010100001011101011100 ;
		12'd 3792 : data_o = 23'b 00010100000111001100101 ;
		12'd 3793 : data_o = 23'b 00010100000010101110000 ;
		12'd 3794 : data_o = 23'b 00010011111110001111011 ;
		12'd 3795 : data_o = 23'b 00010011111001110000111 ;
		12'd 3796 : data_o = 23'b 00010011110101010010100 ;
		12'd 3797 : data_o = 23'b 00010011110000110100010 ;
		12'd 3798 : data_o = 23'b 00010011101100010110001 ;
		12'd 3799 : data_o = 23'b 00010011100111111000001 ;
		12'd 3800 : data_o = 23'b 00010011100011011010001 ;
		12'd 3801 : data_o = 23'b 00010011011110111100011 ;
		12'd 3802 : data_o = 23'b 00010011011010011110101 ;
		12'd 3803 : data_o = 23'b 00010011010110000001000 ;
		12'd 3804 : data_o = 23'b 00010011010001100011100 ;
		12'd 3805 : data_o = 23'b 00010011001101000110001 ;
		12'd 3806 : data_o = 23'b 00010011001000101000110 ;
		12'd 3807 : data_o = 23'b 00010011000100001011101 ;
		12'd 3808 : data_o = 23'b 00010010111111101110100 ;
		12'd 3809 : data_o = 23'b 00010010111011010001101 ;
		12'd 3810 : data_o = 23'b 00010010110110110100110 ;
		12'd 3811 : data_o = 23'b 00010010110010011000000 ;
		12'd 3812 : data_o = 23'b 00010010101101111011011 ;
		12'd 3813 : data_o = 23'b 00010010101001011110111 ;
		12'd 3814 : data_o = 23'b 00010010100101000010011 ;
		12'd 3815 : data_o = 23'b 00010010100000100110001 ;
		12'd 3816 : data_o = 23'b 00010010011100001001111 ;
		12'd 3817 : data_o = 23'b 00010010010111101101110 ;
		12'd 3818 : data_o = 23'b 00010010010011010001110 ;
		12'd 3819 : data_o = 23'b 00010010001110110101111 ;
		12'd 3820 : data_o = 23'b 00010010001010011010001 ;
		12'd 3821 : data_o = 23'b 00010010000101111110100 ;
		12'd 3822 : data_o = 23'b 00010010000001100010111 ;
		12'd 3823 : data_o = 23'b 00010001111101000111100 ;
		12'd 3824 : data_o = 23'b 00010001111000101100001 ;
		12'd 3825 : data_o = 23'b 00010001110100010000111 ;
		12'd 3826 : data_o = 23'b 00010001101111110101110 ;
		12'd 3827 : data_o = 23'b 00010001101011011010110 ;
		12'd 3828 : data_o = 23'b 00010001100110111111110 ;
		12'd 3829 : data_o = 23'b 00010001100010100101000 ;
		12'd 3830 : data_o = 23'b 00010001011110001010010 ;
		12'd 3831 : data_o = 23'b 00010001011001101111101 ;
		12'd 3832 : data_o = 23'b 00010001010101010101010 ;
		12'd 3833 : data_o = 23'b 00010001010000111010111 ;
		12'd 3834 : data_o = 23'b 00010001001100100000100 ;
		12'd 3835 : data_o = 23'b 00010001001000000110011 ;
		12'd 3836 : data_o = 23'b 00010001000011101100010 ;
		12'd 3837 : data_o = 23'b 00010000111111010010011 ;
		12'd 3838 : data_o = 23'b 00010000111010111000100 ;
		12'd 3839 : data_o = 23'b 00010000110110011110110 ;
		12'd 3840 : data_o = 23'b 00010000110010000101001 ;
		12'd 3841 : data_o = 23'b 00010000101101101011101 ;
		12'd 3842 : data_o = 23'b 00010000101001010010001 ;
		12'd 3843 : data_o = 23'b 00010000100100111000111 ;
		12'd 3844 : data_o = 23'b 00010000100000011111101 ;
		12'd 3845 : data_o = 23'b 00010000011100000110100 ;
		12'd 3846 : data_o = 23'b 00010000010111101101100 ;
		12'd 3847 : data_o = 23'b 00010000010011010100101 ;
		12'd 3848 : data_o = 23'b 00010000001110111011111 ;
		12'd 3849 : data_o = 23'b 00010000001010100011010 ;
		12'd 3850 : data_o = 23'b 00010000000110001010101 ;
		12'd 3851 : data_o = 23'b 00010000000001110010001 ;
		12'd 3852 : data_o = 23'b 00001111111101011001110 ;
		12'd 3853 : data_o = 23'b 00001111111001000001100 ;
		12'd 3854 : data_o = 23'b 00001111110100101001011 ;
		12'd 3855 : data_o = 23'b 00001111110000010001011 ;
		12'd 3856 : data_o = 23'b 00001111101011111001011 ;
		12'd 3857 : data_o = 23'b 00001111100111100001101 ;
		12'd 3858 : data_o = 23'b 00001111100011001001111 ;
		12'd 3859 : data_o = 23'b 00001111011110110010010 ;
		12'd 3860 : data_o = 23'b 00001111011010011010110 ;
		12'd 3861 : data_o = 23'b 00001111010110000011010 ;
		12'd 3862 : data_o = 23'b 00001111010001101100000 ;
		12'd 3863 : data_o = 23'b 00001111001101010100110 ;
		12'd 3864 : data_o = 23'b 00001111001000111101110 ;
		12'd 3865 : data_o = 23'b 00001111000100100110110 ;
		12'd 3866 : data_o = 23'b 00001111000000001111111 ;
		12'd 3867 : data_o = 23'b 00001110111011111001000 ;
		12'd 3868 : data_o = 23'b 00001110110111100010011 ;
		12'd 3869 : data_o = 23'b 00001110110011001011110 ;
		12'd 3870 : data_o = 23'b 00001110101110110101011 ;
		12'd 3871 : data_o = 23'b 00001110101010011111000 ;
		12'd 3872 : data_o = 23'b 00001110100110001000110 ;
		12'd 3873 : data_o = 23'b 00001110100001110010101 ;
		12'd 3874 : data_o = 23'b 00001110011101011100100 ;
		12'd 3875 : data_o = 23'b 00001110011001000110101 ;
		12'd 3876 : data_o = 23'b 00001110010100110000110 ;
		12'd 3877 : data_o = 23'b 00001110010000011011000 ;
		12'd 3878 : data_o = 23'b 00001110001100000101011 ;
		12'd 3879 : data_o = 23'b 00001110000111101111111 ;
		12'd 3880 : data_o = 23'b 00001110000011011010100 ;
		12'd 3881 : data_o = 23'b 00001101111111000101001 ;
		12'd 3882 : data_o = 23'b 00001101111010101111111 ;
		12'd 3883 : data_o = 23'b 00001101110110011010110 ;
		12'd 3884 : data_o = 23'b 00001101110010000101110 ;
		12'd 3885 : data_o = 23'b 00001101101101110000111 ;
		12'd 3886 : data_o = 23'b 00001101101001011100001 ;
		12'd 3887 : data_o = 23'b 00001101100101000111011 ;
		12'd 3888 : data_o = 23'b 00001101100000110010111 ;
		12'd 3889 : data_o = 23'b 00001101011100011110011 ;
		12'd 3890 : data_o = 23'b 00001101011000001010000 ;
		12'd 3891 : data_o = 23'b 00001101010011110101110 ;
		12'd 3892 : data_o = 23'b 00001101001111100001100 ;
		12'd 3893 : data_o = 23'b 00001101001011001101100 ;
		12'd 3894 : data_o = 23'b 00001101000110111001100 ;
		12'd 3895 : data_o = 23'b 00001101000010100101101 ;
		12'd 3896 : data_o = 23'b 00001100111110010001111 ;
		12'd 3897 : data_o = 23'b 00001100111001111110010 ;
		12'd 3898 : data_o = 23'b 00001100110101101010110 ;
		12'd 3899 : data_o = 23'b 00001100110001010111010 ;
		12'd 3900 : data_o = 23'b 00001100101101000011111 ;
		12'd 3901 : data_o = 23'b 00001100101000110000101 ;
		12'd 3902 : data_o = 23'b 00001100100100011101100 ;
		12'd 3903 : data_o = 23'b 00001100100000001010100 ;
		12'd 3904 : data_o = 23'b 00001100011011110111101 ;
		12'd 3905 : data_o = 23'b 00001100010111100100110 ;
		12'd 3906 : data_o = 23'b 00001100010011010010000 ;
		12'd 3907 : data_o = 23'b 00001100001110111111011 ;
		12'd 3908 : data_o = 23'b 00001100001010101100111 ;
		12'd 3909 : data_o = 23'b 00001100000110011010100 ;
		12'd 3910 : data_o = 23'b 00001100000010001000001 ;
		12'd 3911 : data_o = 23'b 00001011111101110110000 ;
		12'd 3912 : data_o = 23'b 00001011111001100011111 ;
		12'd 3913 : data_o = 23'b 00001011110101010001111 ;
		12'd 3914 : data_o = 23'b 00001011110000111111111 ;
		12'd 3915 : data_o = 23'b 00001011101100101110001 ;
		12'd 3916 : data_o = 23'b 00001011101000011100011 ;
		12'd 3917 : data_o = 23'b 00001011100100001010111 ;
		12'd 3918 : data_o = 23'b 00001011011111111001011 ;
		12'd 3919 : data_o = 23'b 00001011011011101000000 ;
		12'd 3920 : data_o = 23'b 00001011010111010110101 ;
		12'd 3921 : data_o = 23'b 00001011010011000101100 ;
		12'd 3922 : data_o = 23'b 00001011001110110100011 ;
		12'd 3923 : data_o = 23'b 00001011001010100011011 ;
		12'd 3924 : data_o = 23'b 00001011000110010010100 ;
		12'd 3925 : data_o = 23'b 00001011000010000001110 ;
		12'd 3926 : data_o = 23'b 00001010111101110001001 ;
		12'd 3927 : data_o = 23'b 00001010111001100000100 ;
		12'd 3928 : data_o = 23'b 00001010110101010000001 ;
		12'd 3929 : data_o = 23'b 00001010110000111111110 ;
		12'd 3930 : data_o = 23'b 00001010101100101111011 ;
		12'd 3931 : data_o = 23'b 00001010101000011111010 ;
		12'd 3932 : data_o = 23'b 00001010100100001111010 ;
		12'd 3933 : data_o = 23'b 00001010011111111111010 ;
		12'd 3934 : data_o = 23'b 00001010011011101111011 ;
		12'd 3935 : data_o = 23'b 00001010010111011111101 ;
		12'd 3936 : data_o = 23'b 00001010010011010000000 ;
		12'd 3937 : data_o = 23'b 00001010001111000000011 ;
		12'd 3938 : data_o = 23'b 00001010001010110001000 ;
		12'd 3939 : data_o = 23'b 00001010000110100001101 ;
		12'd 3940 : data_o = 23'b 00001010000010010010011 ;
		12'd 3941 : data_o = 23'b 00001001111110000011010 ;
		12'd 3942 : data_o = 23'b 00001001111001110100001 ;
		12'd 3943 : data_o = 23'b 00001001110101100101010 ;
		12'd 3944 : data_o = 23'b 00001001110001010110011 ;
		12'd 3945 : data_o = 23'b 00001001101101000111101 ;
		12'd 3946 : data_o = 23'b 00001001101000111001000 ;
		12'd 3947 : data_o = 23'b 00001001100100101010011 ;
		12'd 3948 : data_o = 23'b 00001001100000011100000 ;
		12'd 3949 : data_o = 23'b 00001001011100001101101 ;
		12'd 3950 : data_o = 23'b 00001001010111111111011 ;
		12'd 3951 : data_o = 23'b 00001001010011110001010 ;
		12'd 3952 : data_o = 23'b 00001001001111100011010 ;
		12'd 3953 : data_o = 23'b 00001001001011010101010 ;
		12'd 3954 : data_o = 23'b 00001001000111000111100 ;
		12'd 3955 : data_o = 23'b 00001001000010111001110 ;
		12'd 3956 : data_o = 23'b 00001000111110101100001 ;
		12'd 3957 : data_o = 23'b 00001000111010011110100 ;
		12'd 3958 : data_o = 23'b 00001000110110010001001 ;
		12'd 3959 : data_o = 23'b 00001000110010000011110 ;
		12'd 3960 : data_o = 23'b 00001000101101110110100 ;
		12'd 3961 : data_o = 23'b 00001000101001101001011 ;
		12'd 3962 : data_o = 23'b 00001000100101011100011 ;
		12'd 3963 : data_o = 23'b 00001000100001001111011 ;
		12'd 3964 : data_o = 23'b 00001000011101000010101 ;
		12'd 3965 : data_o = 23'b 00001000011000110101111 ;
		12'd 3966 : data_o = 23'b 00001000010100101001010 ;
		12'd 3967 : data_o = 23'b 00001000010000011100110 ;
		12'd 3968 : data_o = 23'b 00001000001100010000010 ;
		12'd 3969 : data_o = 23'b 00001000001000000011111 ;
		12'd 3970 : data_o = 23'b 00001000000011110111101 ;
		12'd 3971 : data_o = 23'b 00000111111111101011100 ;
		12'd 3972 : data_o = 23'b 00000111111011011111100 ;
		12'd 3973 : data_o = 23'b 00000111110111010011101 ;
		12'd 3974 : data_o = 23'b 00000111110011000111110 ;
		12'd 3975 : data_o = 23'b 00000111101110111100000 ;
		12'd 3976 : data_o = 23'b 00000111101010110000011 ;
		12'd 3977 : data_o = 23'b 00000111100110100100111 ;
		12'd 3978 : data_o = 23'b 00000111100010011001011 ;
		12'd 3979 : data_o = 23'b 00000111011110001110000 ;
		12'd 3980 : data_o = 23'b 00000111011010000010110 ;
		12'd 3981 : data_o = 23'b 00000111010101110111101 ;
		12'd 3982 : data_o = 23'b 00000111010001101100101 ;
		12'd 3983 : data_o = 23'b 00000111001101100001101 ;
		12'd 3984 : data_o = 23'b 00000111001001010110111 ;
		12'd 3985 : data_o = 23'b 00000111000101001100001 ;
		12'd 3986 : data_o = 23'b 00000111000001000001100 ;
		12'd 3987 : data_o = 23'b 00000110111100110110111 ;
		12'd 3988 : data_o = 23'b 00000110111000101100100 ;
		12'd 3989 : data_o = 23'b 00000110110100100010001 ;
		12'd 3990 : data_o = 23'b 00000110110000010111111 ;
		12'd 3991 : data_o = 23'b 00000110101100001101110 ;
		12'd 3992 : data_o = 23'b 00000110101000000011101 ;
		12'd 3993 : data_o = 23'b 00000110100011111001110 ;
		12'd 3994 : data_o = 23'b 00000110011111101111111 ;
		12'd 3995 : data_o = 23'b 00000110011011100110001 ;
		12'd 3996 : data_o = 23'b 00000110010111011100011 ;
		12'd 3997 : data_o = 23'b 00000110010011010010111 ;
		12'd 3998 : data_o = 23'b 00000110001111001001011 ;
		12'd 3999 : data_o = 23'b 00000110001011000000000 ;
		12'd 4000 : data_o = 23'b 00000110000110110110110 ;
		12'd 4001 : data_o = 23'b 00000110000010101101101 ;
		12'd 4002 : data_o = 23'b 00000101111110100100100 ;
		12'd 4003 : data_o = 23'b 00000101111010011011101 ;
		12'd 4004 : data_o = 23'b 00000101110110010010110 ;
		12'd 4005 : data_o = 23'b 00000101110010001010000 ;
		12'd 4006 : data_o = 23'b 00000101101110000001010 ;
		12'd 4007 : data_o = 23'b 00000101101001111000101 ;
		12'd 4008 : data_o = 23'b 00000101100101110000010 ;
		12'd 4009 : data_o = 23'b 00000101100001100111111 ;
		12'd 4010 : data_o = 23'b 00000101011101011111100 ;
		12'd 4011 : data_o = 23'b 00000101011001010111011 ;
		12'd 4012 : data_o = 23'b 00000101010101001111010 ;
		12'd 4013 : data_o = 23'b 00000101010001000111010 ;
		12'd 4014 : data_o = 23'b 00000101001100111111011 ;
		12'd 4015 : data_o = 23'b 00000101001000110111101 ;
		12'd 4016 : data_o = 23'b 00000101000100101111111 ;
		12'd 4017 : data_o = 23'b 00000101000000101000010 ;
		12'd 4018 : data_o = 23'b 00000100111100100000110 ;
		12'd 4019 : data_o = 23'b 00000100111000011001011 ;
		12'd 4020 : data_o = 23'b 00000100110100010010001 ;
		12'd 4021 : data_o = 23'b 00000100110000001010111 ;
		12'd 4022 : data_o = 23'b 00000100101100000011110 ;
		12'd 4023 : data_o = 23'b 00000100100111111100110 ;
		12'd 4024 : data_o = 23'b 00000100100011110101111 ;
		12'd 4025 : data_o = 23'b 00000100011111101111000 ;
		12'd 4026 : data_o = 23'b 00000100011011101000010 ;
		12'd 4027 : data_o = 23'b 00000100010111100001101 ;
		12'd 4028 : data_o = 23'b 00000100010011011011001 ;
		12'd 4029 : data_o = 23'b 00000100001111010100101 ;
		12'd 4030 : data_o = 23'b 00000100001011001110011 ;
		12'd 4031 : data_o = 23'b 00000100000111001000001 ;
		12'd 4032 : data_o = 23'b 00000100000011000010000 ;
		12'd 4033 : data_o = 23'b 00000011111110111011111 ;
		12'd 4034 : data_o = 23'b 00000011111010110110000 ;
		12'd 4035 : data_o = 23'b 00000011110110110000001 ;
		12'd 4036 : data_o = 23'b 00000011110010101010011 ;
		12'd 4037 : data_o = 23'b 00000011101110100100110 ;
		12'd 4038 : data_o = 23'b 00000011101010011111001 ;
		12'd 4039 : data_o = 23'b 00000011100110011001101 ;
		12'd 4040 : data_o = 23'b 00000011100010010100010 ;
		12'd 4041 : data_o = 23'b 00000011011110001111000 ;
		12'd 4042 : data_o = 23'b 00000011011010001001111 ;
		12'd 4043 : data_o = 23'b 00000011010110000100110 ;
		12'd 4044 : data_o = 23'b 00000011010001111111110 ;
		12'd 4045 : data_o = 23'b 00000011001101111010111 ;
		12'd 4046 : data_o = 23'b 00000011001001110110001 ;
		12'd 4047 : data_o = 23'b 00000011000101110001011 ;
		12'd 4048 : data_o = 23'b 00000011000001101100110 ;
		12'd 4049 : data_o = 23'b 00000010111101101000010 ;
		12'd 4050 : data_o = 23'b 00000010111001100011111 ;
		12'd 4051 : data_o = 23'b 00000010110101011111100 ;
		12'd 4052 : data_o = 23'b 00000010110001011011011 ;
		12'd 4053 : data_o = 23'b 00000010101101010111010 ;
		12'd 4054 : data_o = 23'b 00000010101001010011010 ;
		12'd 4055 : data_o = 23'b 00000010100101001111010 ;
		12'd 4056 : data_o = 23'b 00000010100001001011011 ;
		12'd 4057 : data_o = 23'b 00000010011101000111110 ;
		12'd 4058 : data_o = 23'b 00000010011001000100000 ;
		12'd 4059 : data_o = 23'b 00000010010101000000100 ;
		12'd 4060 : data_o = 23'b 00000010010000111101000 ;
		12'd 4061 : data_o = 23'b 00000010001100111001110 ;
		12'd 4062 : data_o = 23'b 00000010001000110110011 ;
		12'd 4063 : data_o = 23'b 00000010000100110011010 ;
		12'd 4064 : data_o = 23'b 00000010000000110000010 ;
		12'd 4065 : data_o = 23'b 00000001111100101101010 ;
		12'd 4066 : data_o = 23'b 00000001111000101010011 ;
		12'd 4067 : data_o = 23'b 00000001110100100111100 ;
		12'd 4068 : data_o = 23'b 00000001110000100100111 ;
		12'd 4069 : data_o = 23'b 00000001101100100010010 ;
		12'd 4070 : data_o = 23'b 00000001101000011111110 ;
		12'd 4071 : data_o = 23'b 00000001100100011101011 ;
		12'd 4072 : data_o = 23'b 00000001100000011011000 ;
		12'd 4073 : data_o = 23'b 00000001011100011000111 ;
		12'd 4074 : data_o = 23'b 00000001011000010110110 ;
		12'd 4075 : data_o = 23'b 00000001010100010100101 ;
		12'd 4076 : data_o = 23'b 00000001010000010010110 ;
		12'd 4077 : data_o = 23'b 00000001001100010000111 ;
		12'd 4078 : data_o = 23'b 00000001001000001111001 ;
		12'd 4079 : data_o = 23'b 00000001000100001101100 ;
		12'd 4080 : data_o = 23'b 00000001000000001100000 ;
		12'd 4081 : data_o = 23'b 00000000111100001010100 ;
		12'd 4082 : data_o = 23'b 00000000111000001001001 ;
		12'd 4083 : data_o = 23'b 00000000110100000111111 ;
		12'd 4084 : data_o = 23'b 00000000110000000110110 ;
		12'd 4085 : data_o = 23'b 00000000101100000101101 ;
		12'd 4086 : data_o = 23'b 00000000101000000100101 ;
		12'd 4087 : data_o = 23'b 00000000100100000011110 ;
		12'd 4088 : data_o = 23'b 00000000100000000011000 ;
		12'd 4089 : data_o = 23'b 00000000011100000010010 ;
		12'd 4090 : data_o = 23'b 00000000011000000001101 ;
		12'd 4091 : data_o = 23'b 00000000010100000001001 ;
		12'd 4092 : data_o = 23'b 00000000010000000000110 ;
		12'd 4093 : data_o = 23'b 00000000001100000000011 ;
		12'd 4094 : data_o = 23'b 00000000001000000000001 ;
		12'd 4095 : data_o = 23'b 00000000000100000000000 ;
		default: data_o = 23'd0;
		endcase
	end
endmodule